* NGSPICE file created from spi_slave3.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

.subckt spi_slave3 VGND VPWR clk cs lfsr_seed[0] lfsr_seed[10] lfsr_seed[11] lfsr_seed[12]
+ lfsr_seed[13] lfsr_seed[14] lfsr_seed[15] lfsr_seed[1] lfsr_seed[2] lfsr_seed[3]
+ lfsr_seed[4] lfsr_seed[5] lfsr_seed[6] lfsr_seed[7] lfsr_seed[8] lfsr_seed[9] miso
+ mosi sclk
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_131_ net40 tx_buffer\[3\] _047_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_114_ net29 net8 lfsr_inst.load_seed VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_130_ _050_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_113_ _040_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_8_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold20 _055_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold10 lfsr_inst.lfsr_out\[14\] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
X_112_ net45 net7 lfsr_inst.load_seed VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__mux2_1
Xhold21 lfsr_inst.lfsr_out\[11\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_111_ _039_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold22 _051_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 lfsr_inst.lfsr_out\[9\] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold23 tx_buffer\[4\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
X_110_ net46 net6 lfsr_inst.load_seed VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__mux2_1
Xclkload0 clknet_1_1__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_1
Xhold12 lfsr_inst.lfsr_out\[8\] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold13 _048_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _052_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
X_169_ clknet_1_0__leaf_clk _003_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_15_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold14 tx_buffer\[6\] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_168_ clknet_1_1__leaf_clk _002_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold25 lfsr_inst.lfsr_out\[10\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
X_099_ _033_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold26 lfsr_inst.lfsr_out\[13\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
X_167_ clknet_1_1__leaf_clk _016_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold15 tx_buffer\[1\] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_098_ net23 net15 _066_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_166_ clknet_1_1__leaf_clk _015_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_097_ _032_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold16 tx_buffer\[5\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
X_149_ clknet_1_1__leaf_clk _023_ VGND VGND VPWR VPWR tx_buffer\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold27 lfsr_inst.lfsr_out\[12\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_16_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold17 _053_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_148_ clknet_1_1__leaf_clk _022_ VGND VGND VPWR VPWR tx_buffer\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_7_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_096_ net22 net14 _066_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__mux2_1
X_165_ clknet_1_1__leaf_clk _014_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_16_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_079_ net1 net20 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_164_ clknet_1_1__leaf_clk _013_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[6\] sky130_fd_sc_hd__dfxtp_1
X_095_ _031_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__clkbuf_1
X_078_ _058_ _062_ net1 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__a21oi_1
Xoutput19 net19 VGND VGND VPWR VPWR miso sky130_fd_sc_hd__buf_2
Xhold18 tx_buffer\[2\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_147_ clknet_1_1__leaf_clk _021_ VGND VGND VPWR VPWR tx_buffer\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold19 tx_buffer\[7\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
X_163_ clknet_1_1__leaf_clk _012_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[5\] sky130_fd_sc_hd__dfxtp_1
X_094_ net21 net13 _066_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__mux2_1
X_146_ net18 _020_ VGND VGND VPWR VPWR bit_cnt\[2\] sky130_fd_sc_hd__dfxtp_1
X_077_ bit_cnt\[2\] _059_ _060_ _061_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__a22oi_1
X_129_ lfsr_inst.lfsr_out\[10\] net37 _047_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_162_ clknet_1_0__leaf_clk _011_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_093_ _071_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__clkbuf_1
Xinput1 cs VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_145_ net18 _019_ VGND VGND VPWR VPWR bit_cnt\[1\] sky130_fd_sc_hd__dfxtp_1
X_076_ tx_buffer\[5\] tx_buffer\[4\] bit_cnt\[0\] VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ _049_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 lfsr_seed[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_161_ clknet_1_0__leaf_clk _010_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[3\] sky130_fd_sc_hd__dfxtp_1
X_092_ net27 net12 _066_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_144_ net18 _018_ VGND VGND VPWR VPWR bit_cnt\[0\] sky130_fd_sc_hd__dfxtp_1
X_075_ bit_cnt\[2\] bit_cnt\[1\] VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_11_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_127_ net30 net34 _047_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_143_ net18 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_074_ tx_buffer\[3\] tx_buffer\[2\] tx_buffer\[1\] tx_buffer\[0\] bit_cnt\[0\] bit_cnt\[1\]
+ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_6_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 lfsr_seed[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_160_ clknet_1_0__leaf_clk _009_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[2\] sky130_fd_sc_hd__dfxtp_1
X_091_ _070_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_126_ net32 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_109_ _038_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 lfsr_seed[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_090_ net28 net11 _066_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__mux2_1
X_142_ _056_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
X_073_ bit_cnt\[1\] bit_cnt\[2\] _057_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__or3b_1
X_125_ net31 tx_buffer\[0\] _047_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_108_ net40 net5 lfsr_inst.load_seed VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_141_ net20 _000_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__or2_1
X_072_ tx_buffer\[7\] tx_buffer\[6\] bit_cnt\[0\] VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__mux2_1
Xinput5 lfsr_seed[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_124_ _046_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ _037_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_140_ net39 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 lfsr_seed[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_6_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ bit_cnt\[0\] bit_cnt\[1\] bit_cnt\[2\] seeded VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__or4b_1
X_106_ net44 net4 lfsr_inst.load_seed VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 lfsr_seed[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_122_ bit_cnt\[2\] _045_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__xor2_1
Xinput10 lfsr_seed[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_105_ _036_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 lfsr_seed[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_121_ _044_ _045_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput11 lfsr_seed[3] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_104_ net30 net3 lfsr_inst.load_seed VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput9 lfsr_seed[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_120_ bit_cnt\[1\] _042_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 lfsr_seed[4] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_103_ _035_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__clkbuf_1
Xhold1 seeded VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_102_ net31 net17 _066_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__mux2_1
Xinput13 lfsr_seed[5] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_13_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold2 lfsr_inst.lfsr_out\[4\] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 lfsr_seed[6] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_101_ _034_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 lfsr_inst.lfsr_out\[5\] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 lfsr_seed[7] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_100_ net25 net16 _066_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 lfsr_inst.lfsr_out\[6\] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 lfsr_seed[8] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_159_ clknet_1_0__leaf_clk _008_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold5 lfsr_inst.lfsr_out\[1\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_17_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 lfsr_seed[9] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_158_ clknet_1_0__leaf_clk _001_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_5_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ _069_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__clkbuf_1
Xhold6 lfsr_inst.lfsr_out\[7\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput18 sclk VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
X_157_ _017_ _030_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_1
X_088_ net24 net10 _066_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold7 lfsr_inst.lfsr_out\[0\] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_173_ clknet_1_0__leaf_clk _007_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_156_ clknet_1_1__leaf_clk _029_ VGND VGND VPWR VPWR seeded sky130_fd_sc_hd__dfxtp_1
X_087_ _068_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__clkbuf_1
Xhold8 lfsr_inst.lfsr_out\[3\] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
X_139_ lfsr_inst.lfsr_out\[15\] net38 _047_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_155_ clknet_1_1__leaf_clk _000_ VGND VGND VPWR VPWR lfsr_inst.load_seed sky130_fd_sc_hd__dfxtp_2
X_172_ clknet_1_0__leaf_clk _006_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[14\] sky130_fd_sc_hd__dfxtp_1
X_086_ net26 net9 _066_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__mux2_1
X_138_ _054_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold9 lfsr_inst.lfsr_out\[2\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_171_ clknet_1_0__leaf_clk _005_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[13\] sky130_fd_sc_hd__dfxtp_1
X_154_ clknet_1_0__leaf_clk _028_ VGND VGND VPWR VPWR tx_buffer\[7\] sky130_fd_sc_hd__dfxtp_1
X_085_ _067_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
X_137_ net29 net33 _047_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ clknet_1_0__leaf_clk _004_ VGND VGND VPWR VPWR lfsr_inst.lfsr_out\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_153_ clknet_1_0__leaf_clk _027_ VGND VGND VPWR VPWR tx_buffer\[6\] sky130_fd_sc_hd__dfxtp_1
X_136_ net36 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_084_ _065_ net2 _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_119_ bit_cnt\[1\] _042_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ clknet_1_0__leaf_clk _026_ VGND VGND VPWR VPWR tx_buffer\[5\] sky130_fd_sc_hd__dfxtp_1
X_083_ lfsr_inst.load_seed VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__clkbuf_4
X_118_ _042_ _043_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__nor2_1
X_135_ lfsr_inst.lfsr_out\[13\] net35 _047_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_151_ clknet_1_0__leaf_clk _025_ VGND VGND VPWR VPWR tx_buffer\[4\] sky130_fd_sc_hd__dfxtp_1
X_134_ net43 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
X_082_ _063_ _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ bit_cnt\[0\] net1 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__and2b_1
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_081_ lfsr_inst.lfsr_out\[15\] lfsr_inst.lfsr_out\[13\] VGND VGND VPWR VPWR _064_
+ sky130_fd_sc_hd__xor2_1
X_150_ clknet_1_1__leaf_clk _024_ VGND VGND VPWR VPWR tx_buffer\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_133_ lfsr_inst.lfsr_out\[12\] net42 _047_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_116_ net1 bit_cnt\[0\] VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_132_ net41 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__clkbuf_1
X_080_ lfsr_inst.lfsr_out\[12\] lfsr_inst.lfsr_out\[10\] VGND VGND VPWR VPWR _063_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_115_ _041_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

