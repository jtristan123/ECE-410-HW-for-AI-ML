magic
tech sky130A
magscale 1 2
timestamp 1749864851
<< checkpaint >>
rect -3932 -3932 16054 18198
<< viali >>
rect 4813 11713 4847 11747
rect 5273 11713 5307 11747
rect 7849 11713 7883 11747
rect 5089 11577 5123 11611
rect 4629 11509 4663 11543
rect 8033 11509 8067 11543
rect 5365 11305 5399 11339
rect 4537 11237 4571 11271
rect 3985 11169 4019 11203
rect 5917 11169 5951 11203
rect 7205 11169 7239 11203
rect 2421 11101 2455 11135
rect 4169 11101 4203 11135
rect 4629 11101 4663 11135
rect 5181 11101 5215 11135
rect 6101 11101 6135 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 7757 11101 7791 11135
rect 7941 11101 7975 11135
rect 8125 11101 8159 11135
rect 4077 11033 4111 11067
rect 6561 11033 6595 11067
rect 8033 11033 8067 11067
rect 2237 10965 2271 10999
rect 6285 10965 6319 10999
rect 3341 10761 3375 10795
rect 4997 10761 5031 10795
rect 5825 10761 5859 10795
rect 7757 10761 7791 10795
rect 3884 10693 3918 10727
rect 5089 10693 5123 10727
rect 6193 10693 6227 10727
rect 6622 10693 6656 10727
rect 8962 10693 8996 10727
rect 1409 10625 1443 10659
rect 1961 10625 1995 10659
rect 2228 10625 2262 10659
rect 6009 10625 6043 10659
rect 3617 10557 3651 10591
rect 5641 10557 5675 10591
rect 6377 10557 6411 10591
rect 9229 10557 9263 10591
rect 1593 10421 1627 10455
rect 7849 10421 7883 10455
rect 2329 10217 2363 10251
rect 5181 10217 5215 10251
rect 7481 10217 7515 10251
rect 8125 10217 8159 10251
rect 8217 10217 8251 10251
rect 10425 10217 10459 10251
rect 7941 10149 7975 10183
rect 8401 10149 8435 10183
rect 2789 10081 2823 10115
rect 2973 10081 3007 10115
rect 3801 10081 3835 10115
rect 8677 10081 8711 10115
rect 10333 10081 10367 10115
rect 4068 10013 4102 10047
rect 6837 10013 6871 10047
rect 7113 10013 7147 10047
rect 7297 10013 7331 10047
rect 7573 10013 7607 10047
rect 10609 10013 10643 10047
rect 6570 9945 6604 9979
rect 7665 9945 7699 9979
rect 10066 9945 10100 9979
rect 2697 9877 2731 9911
rect 5457 9877 5491 9911
rect 6929 9877 6963 9911
rect 8953 9877 8987 9911
rect 5273 9673 5307 9707
rect 4077 9605 4111 9639
rect 1685 9537 1719 9571
rect 1952 9537 1986 9571
rect 3525 9537 3559 9571
rect 4169 9537 4203 9571
rect 5181 9537 5215 9571
rect 6929 9537 6963 9571
rect 7021 9537 7055 9571
rect 7389 9537 7423 9571
rect 7941 9537 7975 9571
rect 8033 9537 8067 9571
rect 8493 9537 8527 9571
rect 10066 9537 10100 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 3433 9469 3467 9503
rect 3985 9469 4019 9503
rect 5089 9469 5123 9503
rect 8217 9469 8251 9503
rect 8401 9469 8435 9503
rect 8861 9469 8895 9503
rect 4537 9401 4571 9435
rect 5641 9401 5675 9435
rect 8953 9401 8987 9435
rect 3065 9333 3099 9367
rect 3157 9333 3191 9367
rect 6745 9333 6779 9367
rect 7297 9333 7331 9367
rect 7573 9333 7607 9367
rect 10517 9333 10551 9367
rect 1961 9129 1995 9163
rect 3617 9129 3651 9163
rect 8493 9129 8527 9163
rect 4813 9061 4847 9095
rect 7297 9061 7331 9095
rect 3065 8993 3099 9027
rect 4261 8993 4295 9027
rect 6285 8993 6319 9027
rect 8125 8993 8159 9027
rect 9045 8993 9079 9027
rect 2145 8925 2179 8959
rect 5641 8925 5675 8959
rect 7481 8925 7515 8959
rect 7573 8925 7607 8959
rect 8033 8925 8067 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 8493 8925 8527 8959
rect 9301 8925 9335 8959
rect 4353 8857 4387 8891
rect 4997 8857 5031 8891
rect 7297 8857 7331 8891
rect 4445 8789 4479 8823
rect 5733 8789 5767 8823
rect 10425 8789 10459 8823
rect 2237 8585 2271 8619
rect 5365 8585 5399 8619
rect 5825 8585 5859 8619
rect 6193 8585 6227 8619
rect 10517 8585 10551 8619
rect 7389 8517 7423 8551
rect 7941 8517 7975 8551
rect 8217 8517 8251 8551
rect 1409 8449 1443 8483
rect 2605 8449 2639 8483
rect 3065 8449 3099 8483
rect 4252 8449 4286 8483
rect 8125 8449 8159 8483
rect 8345 8449 8379 8483
rect 10333 8449 10367 8483
rect 2697 8381 2731 8415
rect 2789 8381 2823 8415
rect 3617 8381 3651 8415
rect 3985 8381 4019 8415
rect 5641 8381 5675 8415
rect 5733 8381 5767 8415
rect 7849 8381 7883 8415
rect 1593 8313 1627 8347
rect 7665 8313 7699 8347
rect 7941 8313 7975 8347
rect 3065 8041 3099 8075
rect 3985 8041 4019 8075
rect 5641 8041 5675 8075
rect 1685 7905 1719 7939
rect 1409 7837 1443 7871
rect 3433 7837 3467 7871
rect 3801 7837 3835 7871
rect 4261 7837 4295 7871
rect 6745 7837 6779 7871
rect 8125 7837 8159 7871
rect 9965 7837 9999 7871
rect 1952 7769 1986 7803
rect 4506 7769 4540 7803
rect 1593 7701 1627 7735
rect 3617 7701 3651 7735
rect 6561 7701 6595 7735
rect 8677 7701 8711 7735
rect 10517 7701 10551 7735
rect 1961 7497 1995 7531
rect 2237 7497 2271 7531
rect 2697 7497 2731 7531
rect 7757 7497 7791 7531
rect 9781 7497 9815 7531
rect 1409 7361 1443 7395
rect 2145 7361 2179 7395
rect 2605 7361 2639 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 6644 7361 6678 7395
rect 7941 7361 7975 7395
rect 9137 7361 9171 7395
rect 9873 7361 9907 7395
rect 2789 7293 2823 7327
rect 6377 7293 6411 7327
rect 8125 7293 8159 7327
rect 8861 7293 8895 7327
rect 8978 7293 9012 7327
rect 8585 7225 8619 7259
rect 1593 7157 1627 7191
rect 3893 7157 3927 7191
rect 5273 7157 5307 7191
rect 10517 7157 10551 7191
rect 5181 6953 5215 6987
rect 7849 6953 7883 6987
rect 3341 6817 3375 6851
rect 4445 6817 4479 6851
rect 4629 6817 4663 6851
rect 8309 6817 8343 6851
rect 8401 6817 8435 6851
rect 1593 6749 1627 6783
rect 3433 6749 3467 6783
rect 5733 6749 5767 6783
rect 6009 6749 6043 6783
rect 10333 6749 10367 6783
rect 10609 6749 10643 6783
rect 1860 6681 1894 6715
rect 8217 6681 8251 6715
rect 10088 6681 10122 6715
rect 2973 6613 3007 6647
rect 3065 6613 3099 6647
rect 4721 6613 4755 6647
rect 5089 6613 5123 6647
rect 7297 6613 7331 6647
rect 8953 6613 8987 6647
rect 10425 6613 10459 6647
rect 1869 6409 1903 6443
rect 2145 6409 2179 6443
rect 2605 6409 2639 6443
rect 2973 6409 3007 6443
rect 3709 6409 3743 6443
rect 6193 6409 6227 6443
rect 9689 6409 9723 6443
rect 2513 6341 2547 6375
rect 7849 6341 7883 6375
rect 1409 6273 1443 6307
rect 2053 6273 2087 6307
rect 3617 6273 3651 6307
rect 4077 6273 4111 6307
rect 4701 6273 4735 6307
rect 6009 6273 6043 6307
rect 6377 6273 6411 6307
rect 6633 6273 6667 6307
rect 10609 6273 10643 6307
rect 2697 6205 2731 6239
rect 3985 6205 4019 6239
rect 4445 6205 4479 6239
rect 9597 6205 9631 6239
rect 10241 6205 10275 6239
rect 5825 6137 5859 6171
rect 1593 6069 1627 6103
rect 7757 6069 7791 6103
rect 10425 6069 10459 6103
rect 7205 5865 7239 5899
rect 8769 5865 8803 5899
rect 8953 5865 8987 5899
rect 3617 5797 3651 5831
rect 3065 5729 3099 5763
rect 4905 5729 4939 5763
rect 5089 5729 5123 5763
rect 6745 5729 6779 5763
rect 7849 5729 7883 5763
rect 8125 5729 8159 5763
rect 8309 5729 8343 5763
rect 1409 5661 1443 5695
rect 3249 5661 3283 5695
rect 3893 5661 3927 5695
rect 10333 5661 10367 5695
rect 4813 5593 4847 5627
rect 6478 5593 6512 5627
rect 8401 5593 8435 5627
rect 10088 5593 10122 5627
rect 1593 5525 1627 5559
rect 3157 5525 3191 5559
rect 3985 5525 4019 5559
rect 4445 5525 4479 5559
rect 5365 5525 5399 5559
rect 6929 5525 6963 5559
rect 7573 5525 7607 5559
rect 7665 5525 7699 5559
rect 3985 5321 4019 5355
rect 4721 5321 4755 5355
rect 5549 5321 5583 5355
rect 6377 5321 6411 5355
rect 9321 5321 9355 5355
rect 9781 5321 9815 5355
rect 2044 5253 2078 5287
rect 1409 5185 1443 5219
rect 4169 5185 4203 5219
rect 4537 5185 4571 5219
rect 6193 5185 6227 5219
rect 6561 5185 6595 5219
rect 8053 5185 8087 5219
rect 8309 5185 8343 5219
rect 9413 5185 9447 5219
rect 10241 5185 10275 5219
rect 1777 5117 1811 5151
rect 3801 5117 3835 5151
rect 9137 5117 9171 5151
rect 10333 5117 10367 5151
rect 10425 5117 10459 5151
rect 3157 5049 3191 5083
rect 9873 5049 9907 5083
rect 1593 4981 1627 5015
rect 3249 4981 3283 5015
rect 6929 4981 6963 5015
rect 6745 4777 6779 4811
rect 6837 4777 6871 4811
rect 7757 4777 7791 4811
rect 8493 4777 8527 4811
rect 10425 4777 10459 4811
rect 2513 4709 2547 4743
rect 5089 4709 5123 4743
rect 2973 4641 3007 4675
rect 3157 4641 3191 4675
rect 6101 4641 6135 4675
rect 7389 4641 7423 4675
rect 8401 4641 8435 4675
rect 8953 4641 8987 4675
rect 2329 4573 2363 4607
rect 2881 4573 2915 4607
rect 4353 4573 4387 4607
rect 4629 4573 4663 4607
rect 4905 4573 4939 4607
rect 5825 4573 5859 4607
rect 6377 4573 6411 4607
rect 8677 4573 8711 4607
rect 10609 4573 10643 4607
rect 9220 4505 9254 4539
rect 2145 4437 2179 4471
rect 3801 4437 3835 4471
rect 4813 4437 4847 4471
rect 5181 4437 5215 4471
rect 6285 4437 6319 4471
rect 10333 4437 10367 4471
rect 4721 4233 4755 4267
rect 5089 4233 5123 4267
rect 6377 4233 6411 4267
rect 9597 4233 9631 4267
rect 9873 4233 9907 4267
rect 2044 4165 2078 4199
rect 9137 4165 9171 4199
rect 3525 4097 3559 4131
rect 6193 4097 6227 4131
rect 6745 4097 6779 4131
rect 8309 4097 8343 4131
rect 9781 4097 9815 4131
rect 10425 4097 10459 4131
rect 1777 4029 1811 4063
rect 3801 4029 3835 4063
rect 5181 4029 5215 4063
rect 5365 4029 5399 4063
rect 5641 4029 5675 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7757 4029 7791 4063
rect 8125 4029 8159 4063
rect 8217 4029 8251 4063
rect 8861 4029 8895 4063
rect 9045 4029 9079 4063
rect 3157 3961 3191 3995
rect 9505 3961 9539 3995
rect 3709 3893 3743 3927
rect 4445 3893 4479 3927
rect 7205 3893 7239 3927
rect 8677 3893 8711 3927
rect 3617 3689 3651 3723
rect 5181 3689 5215 3723
rect 6837 3689 6871 3723
rect 8953 3689 8987 3723
rect 9689 3689 9723 3723
rect 10425 3689 10459 3723
rect 8309 3621 8343 3655
rect 9505 3553 9539 3587
rect 1961 3485 1995 3519
rect 2237 3485 2271 3519
rect 3801 3485 3835 3519
rect 5457 3485 5491 3519
rect 6929 3485 6963 3519
rect 8585 3485 8619 3519
rect 10241 3485 10275 3519
rect 10609 3485 10643 3519
rect 2482 3417 2516 3451
rect 4046 3417 4080 3451
rect 5724 3417 5758 3451
rect 7196 3417 7230 3451
rect 2145 3349 2179 3383
rect 8401 3349 8435 3383
rect 2697 3145 2731 3179
rect 3065 3145 3099 3179
rect 3617 3145 3651 3179
rect 3985 3145 4019 3179
rect 6193 3145 6227 3179
rect 7205 3145 7239 3179
rect 7573 3145 7607 3179
rect 7665 3145 7699 3179
rect 9413 3145 9447 3179
rect 4077 3077 4111 3111
rect 5080 3077 5114 3111
rect 4813 3009 4847 3043
rect 7849 3009 7883 3043
rect 8033 3009 8067 3043
rect 8300 3009 8334 3043
rect 3157 2941 3191 2975
rect 3341 2941 3375 2975
rect 4261 2941 4295 2975
rect 7021 2941 7055 2975
rect 7113 2941 7147 2975
rect 3341 2601 3375 2635
rect 4169 2601 4203 2635
rect 5273 2601 5307 2635
rect 6101 2601 6135 2635
rect 6561 2601 6595 2635
rect 7205 2601 7239 2635
rect 8493 2601 8527 2635
rect 3525 2397 3559 2431
rect 3985 2397 4019 2431
rect 5457 2397 5491 2431
rect 5917 2397 5951 2431
rect 6745 2397 6779 2431
rect 7389 2397 7423 2431
rect 8677 2397 8711 2431
<< metal1 >>
rect 1104 11994 10948 12016
rect 1104 11942 2840 11994
rect 2892 11942 2904 11994
rect 2956 11942 2968 11994
rect 3020 11942 3032 11994
rect 3084 11942 3096 11994
rect 3148 11942 5301 11994
rect 5353 11942 5365 11994
rect 5417 11942 5429 11994
rect 5481 11942 5493 11994
rect 5545 11942 5557 11994
rect 5609 11942 7762 11994
rect 7814 11942 7826 11994
rect 7878 11942 7890 11994
rect 7942 11942 7954 11994
rect 8006 11942 8018 11994
rect 8070 11942 10223 11994
rect 10275 11942 10287 11994
rect 10339 11942 10351 11994
rect 10403 11942 10415 11994
rect 10467 11942 10479 11994
rect 10531 11942 10948 11994
rect 1104 11920 10948 11942
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 5166 11744 5172 11756
rect 4847 11716 5172 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 5166 11704 5172 11716
rect 5224 11704 5230 11756
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 4522 11636 4528 11688
rect 4580 11676 4586 11688
rect 5276 11676 5304 11707
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 7708 11716 7849 11744
rect 7708 11704 7714 11716
rect 7837 11713 7849 11716
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 4580 11648 5304 11676
rect 4580 11636 4586 11648
rect 4154 11568 4160 11620
rect 4212 11608 4218 11620
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4212 11580 5089 11608
rect 4212 11568 4218 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5077 11571 5135 11577
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4396 11512 4629 11540
rect 4396 11500 4402 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7616 11512 8033 11540
rect 7616 11500 7622 11512
rect 8021 11509 8033 11512
rect 8067 11509 8079 11543
rect 8021 11503 8079 11509
rect 1104 11450 10948 11472
rect 1104 11398 2180 11450
rect 2232 11398 2244 11450
rect 2296 11398 2308 11450
rect 2360 11398 2372 11450
rect 2424 11398 2436 11450
rect 2488 11398 4641 11450
rect 4693 11398 4705 11450
rect 4757 11398 4769 11450
rect 4821 11398 4833 11450
rect 4885 11398 4897 11450
rect 4949 11398 7102 11450
rect 7154 11398 7166 11450
rect 7218 11398 7230 11450
rect 7282 11398 7294 11450
rect 7346 11398 7358 11450
rect 7410 11398 9563 11450
rect 9615 11398 9627 11450
rect 9679 11398 9691 11450
rect 9743 11398 9755 11450
rect 9807 11398 9819 11450
rect 9871 11398 10948 11450
rect 1104 11376 10948 11398
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 5353 11339 5411 11345
rect 5353 11336 5365 11339
rect 5224 11308 5365 11336
rect 5224 11296 5230 11308
rect 5353 11305 5365 11308
rect 5399 11305 5411 11339
rect 5353 11299 5411 11305
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11268 4583 11271
rect 4571 11240 5948 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 3973 11203 4031 11209
rect 3973 11169 3985 11203
rect 4019 11200 4031 11203
rect 4430 11200 4436 11212
rect 4019 11172 4436 11200
rect 4019 11169 4031 11172
rect 3973 11163 4031 11169
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 5920 11209 5948 11240
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11169 5963 11203
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 5905 11163 5963 11169
rect 6472 11172 7205 11200
rect 6472 11144 6500 11172
rect 7193 11169 7205 11172
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2498 11132 2504 11144
rect 2455 11104 2504 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2498 11092 2504 11104
rect 2556 11092 2562 11144
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 4157 11135 4215 11141
rect 4157 11132 4169 11135
rect 3384 11104 4169 11132
rect 3384 11092 3390 11104
rect 4157 11101 4169 11104
rect 4203 11101 4215 11135
rect 4157 11095 4215 11101
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4304 11104 4629 11132
rect 4304 11092 4310 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 5166 11092 5172 11144
rect 5224 11092 5230 11144
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 6454 11092 6460 11144
rect 6512 11092 6518 11144
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 7558 11132 7564 11144
rect 6687 11104 7564 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7745 11135 7803 11141
rect 7745 11132 7757 11135
rect 7708 11104 7757 11132
rect 7708 11092 7714 11104
rect 7745 11101 7757 11104
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 4890 11064 4896 11076
rect 4111 11036 4896 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 6178 11024 6184 11076
rect 6236 11064 6242 11076
rect 6549 11067 6607 11073
rect 6549 11064 6561 11067
rect 6236 11036 6561 11064
rect 6236 11024 6242 11036
rect 6549 11033 6561 11036
rect 6595 11033 6607 11067
rect 6549 11027 6607 11033
rect 2222 10956 2228 11008
rect 2280 10956 2286 11008
rect 6270 10956 6276 11008
rect 6328 10956 6334 11008
rect 7944 10996 7972 11095
rect 8110 11092 8116 11144
rect 8168 11092 8174 11144
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 8938 11064 8944 11076
rect 8067 11036 8944 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 8202 10996 8208 11008
rect 7944 10968 8208 10996
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 1104 10906 10948 10928
rect 1104 10854 2840 10906
rect 2892 10854 2904 10906
rect 2956 10854 2968 10906
rect 3020 10854 3032 10906
rect 3084 10854 3096 10906
rect 3148 10854 5301 10906
rect 5353 10854 5365 10906
rect 5417 10854 5429 10906
rect 5481 10854 5493 10906
rect 5545 10854 5557 10906
rect 5609 10854 7762 10906
rect 7814 10854 7826 10906
rect 7878 10854 7890 10906
rect 7942 10854 7954 10906
rect 8006 10854 8018 10906
rect 8070 10854 10223 10906
rect 10275 10854 10287 10906
rect 10339 10854 10351 10906
rect 10403 10854 10415 10906
rect 10467 10854 10479 10906
rect 10531 10854 10948 10906
rect 1104 10832 10948 10854
rect 3326 10752 3332 10804
rect 3384 10752 3390 10804
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 5166 10792 5172 10804
rect 5031 10764 5172 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 6086 10792 6092 10804
rect 5859 10764 6092 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 7708 10764 7757 10792
rect 7708 10752 7714 10764
rect 7745 10761 7757 10764
rect 7791 10761 7803 10795
rect 7745 10755 7803 10761
rect 3872 10727 3930 10733
rect 1964 10696 3648 10724
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 900 10628 1409 10656
rect 900 10616 906 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 1670 10616 1676 10668
rect 1728 10656 1734 10668
rect 1964 10665 1992 10696
rect 2222 10665 2228 10668
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1728 10628 1961 10656
rect 1728 10616 1734 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 2216 10656 2228 10665
rect 2183 10628 2228 10656
rect 1949 10619 2007 10625
rect 2216 10619 2228 10628
rect 2222 10616 2228 10619
rect 2280 10616 2286 10668
rect 3620 10600 3648 10696
rect 3872 10693 3884 10727
rect 3918 10724 3930 10727
rect 4154 10724 4160 10736
rect 3918 10696 4160 10724
rect 3918 10693 3930 10696
rect 3872 10687 3930 10693
rect 4154 10684 4160 10696
rect 4212 10684 4218 10736
rect 4890 10684 4896 10736
rect 4948 10724 4954 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 4948 10696 5089 10724
rect 4948 10684 4954 10696
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 6178 10684 6184 10736
rect 6236 10684 6242 10736
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 6610 10727 6668 10733
rect 6610 10724 6622 10727
rect 6328 10696 6622 10724
rect 6328 10684 6334 10696
rect 6610 10693 6622 10696
rect 6656 10693 6668 10727
rect 6610 10687 6668 10693
rect 8938 10684 8944 10736
rect 8996 10733 9002 10736
rect 8996 10724 9008 10733
rect 8996 10696 9041 10724
rect 8996 10687 9008 10696
rect 8996 10684 9002 10687
rect 5997 10659 6055 10665
rect 5997 10625 6009 10659
rect 6043 10656 6055 10659
rect 6454 10656 6460 10668
rect 6043 10628 6460 10656
rect 6043 10625 6055 10628
rect 5997 10619 6055 10625
rect 6454 10616 6460 10628
rect 6512 10616 6518 10668
rect 3602 10548 3608 10600
rect 3660 10548 3666 10600
rect 5166 10548 5172 10600
rect 5224 10588 5230 10600
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 5224 10560 5641 10588
rect 5224 10548 5230 10560
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 6362 10548 6368 10600
rect 6420 10548 6426 10600
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10588 9275 10591
rect 10410 10588 10416 10600
rect 9263 10560 10416 10588
rect 9263 10557 9275 10560
rect 9217 10551 9275 10557
rect 10410 10548 10416 10560
rect 10468 10548 10474 10600
rect 1578 10412 1584 10464
rect 1636 10412 1642 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7834 10452 7840 10464
rect 7064 10424 7840 10452
rect 7064 10412 7070 10424
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 1104 10362 10948 10384
rect 1104 10310 2180 10362
rect 2232 10310 2244 10362
rect 2296 10310 2308 10362
rect 2360 10310 2372 10362
rect 2424 10310 2436 10362
rect 2488 10310 4641 10362
rect 4693 10310 4705 10362
rect 4757 10310 4769 10362
rect 4821 10310 4833 10362
rect 4885 10310 4897 10362
rect 4949 10310 7102 10362
rect 7154 10310 7166 10362
rect 7218 10310 7230 10362
rect 7282 10310 7294 10362
rect 7346 10310 7358 10362
rect 7410 10310 9563 10362
rect 9615 10310 9627 10362
rect 9679 10310 9691 10362
rect 9743 10310 9755 10362
rect 9807 10310 9819 10362
rect 9871 10310 10948 10362
rect 1104 10288 10948 10310
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2498 10248 2504 10260
rect 2363 10220 2504 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 5166 10208 5172 10260
rect 5224 10208 5230 10260
rect 7469 10251 7527 10257
rect 7469 10217 7481 10251
rect 7515 10217 7527 10251
rect 7469 10211 7527 10217
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 1636 10084 2789 10112
rect 1636 10072 1642 10084
rect 2777 10081 2789 10084
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3007 10084 3372 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 2682 10004 2688 10056
rect 2740 10044 2746 10056
rect 2976 10044 3004 10075
rect 2740 10016 3004 10044
rect 2740 10004 2746 10016
rect 3344 9976 3372 10084
rect 3602 10072 3608 10124
rect 3660 10112 3666 10124
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 3660 10084 3801 10112
rect 3660 10072 3666 10084
rect 3789 10081 3801 10084
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 4056 10047 4114 10053
rect 4056 10013 4068 10047
rect 4102 10044 4114 10047
rect 4338 10044 4344 10056
rect 4102 10016 4344 10044
rect 4102 10013 4114 10016
rect 4056 10007 4114 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6380 10016 6837 10044
rect 6380 9988 6408 10016
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 7064 10016 7113 10044
rect 7064 10004 7070 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 7282 10004 7288 10056
rect 7340 10004 7346 10056
rect 3344 9948 5488 9976
rect 2685 9911 2743 9917
rect 2685 9877 2697 9911
rect 2731 9908 2743 9911
rect 3602 9908 3608 9920
rect 2731 9880 3608 9908
rect 2731 9877 2743 9880
rect 2685 9871 2743 9877
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 5460 9917 5488 9948
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 6558 9979 6616 9985
rect 6558 9976 6570 9979
rect 6472 9948 6570 9976
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9877 5503 9911
rect 5445 9871 5503 9877
rect 6178 9868 6184 9920
rect 6236 9908 6242 9920
rect 6472 9908 6500 9948
rect 6558 9945 6570 9948
rect 6604 9945 6616 9979
rect 7484 9976 7512 10211
rect 8110 10208 8116 10260
rect 8168 10208 8174 10260
rect 8202 10208 8208 10260
rect 8260 10208 8266 10260
rect 10410 10208 10416 10260
rect 10468 10208 10474 10260
rect 7742 10140 7748 10192
rect 7800 10180 7806 10192
rect 7929 10183 7987 10189
rect 7929 10180 7941 10183
rect 7800 10152 7941 10180
rect 7800 10140 7806 10152
rect 7929 10149 7941 10152
rect 7975 10149 7987 10183
rect 7929 10143 7987 10149
rect 8389 10183 8447 10189
rect 8389 10149 8401 10183
rect 8435 10180 8447 10183
rect 8570 10180 8576 10192
rect 8435 10152 8576 10180
rect 8435 10149 8447 10152
rect 8389 10143 8447 10149
rect 7650 10112 7656 10124
rect 7576 10084 7656 10112
rect 7576 10053 7604 10084
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 7944 10112 7972 10143
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 8665 10115 8723 10121
rect 8665 10112 8677 10115
rect 7944 10084 8677 10112
rect 8665 10081 8677 10084
rect 8711 10081 8723 10115
rect 8665 10075 8723 10081
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 10428 10112 10456 10208
rect 10686 10112 10692 10124
rect 10367 10084 10692 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 10686 10072 10692 10084
rect 10744 10072 10750 10124
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 7653 9979 7711 9985
rect 7484 9948 7604 9976
rect 6558 9939 6616 9945
rect 6236 9880 6500 9908
rect 6236 9868 6242 9880
rect 6914 9868 6920 9920
rect 6972 9868 6978 9920
rect 7576 9908 7604 9948
rect 7653 9945 7665 9979
rect 7699 9976 7711 9979
rect 7834 9976 7840 9988
rect 7699 9948 7840 9976
rect 7699 9945 7711 9948
rect 7653 9939 7711 9945
rect 7834 9936 7840 9948
rect 7892 9976 7898 9988
rect 8570 9976 8576 9988
rect 7892 9948 8576 9976
rect 7892 9936 7898 9948
rect 8570 9936 8576 9948
rect 8628 9936 8634 9988
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 10054 9979 10112 9985
rect 10054 9976 10066 9979
rect 9272 9948 10066 9976
rect 9272 9936 9278 9948
rect 10054 9945 10066 9948
rect 10100 9945 10112 9979
rect 10054 9939 10112 9945
rect 8294 9908 8300 9920
rect 7576 9880 8300 9908
rect 8294 9868 8300 9880
rect 8352 9908 8358 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8352 9880 8953 9908
rect 8352 9868 8358 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 1104 9818 10948 9840
rect 1104 9766 2840 9818
rect 2892 9766 2904 9818
rect 2956 9766 2968 9818
rect 3020 9766 3032 9818
rect 3084 9766 3096 9818
rect 3148 9766 5301 9818
rect 5353 9766 5365 9818
rect 5417 9766 5429 9818
rect 5481 9766 5493 9818
rect 5545 9766 5557 9818
rect 5609 9766 7762 9818
rect 7814 9766 7826 9818
rect 7878 9766 7890 9818
rect 7942 9766 7954 9818
rect 8006 9766 8018 9818
rect 8070 9766 10223 9818
rect 10275 9766 10287 9818
rect 10339 9766 10351 9818
rect 10403 9766 10415 9818
rect 10467 9766 10479 9818
rect 10531 9766 10948 9818
rect 1104 9744 10948 9766
rect 5166 9664 5172 9716
rect 5224 9704 5230 9716
rect 5261 9707 5319 9713
rect 5261 9704 5273 9707
rect 5224 9676 5273 9704
rect 5224 9664 5230 9676
rect 5261 9673 5273 9676
rect 5307 9673 5319 9707
rect 8294 9704 8300 9716
rect 5261 9667 5319 9673
rect 8036 9676 8300 9704
rect 4065 9639 4123 9645
rect 4065 9605 4077 9639
rect 4111 9636 4123 9639
rect 4246 9636 4252 9648
rect 4111 9608 4252 9636
rect 4111 9605 4123 9608
rect 4065 9599 4123 9605
rect 4246 9596 4252 9608
rect 4304 9596 4310 9648
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 8036 9636 8064 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 5132 9608 5212 9636
rect 5132 9596 5138 9608
rect 1670 9528 1676 9580
rect 1728 9528 1734 9580
rect 1946 9577 1952 9580
rect 1940 9531 1952 9577
rect 1946 9528 1952 9531
rect 2004 9528 2010 9580
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 3384 9540 3525 9568
rect 3384 9528 3390 9540
rect 3513 9537 3525 9540
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 5184 9577 5212 9608
rect 7944 9608 8064 9636
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 3660 9540 4169 9568
rect 3660 9528 3666 9540
rect 4157 9537 4169 9540
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7944 9577 7972 9608
rect 8202 9596 8208 9648
rect 8260 9596 8266 9648
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9568 7435 9571
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7423 9540 7941 9568
rect 7423 9537 7435 9540
rect 7377 9531 7435 9537
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 7929 9531 7987 9537
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8220 9568 8248 9596
rect 8067 9540 8248 9568
rect 8481 9571 8539 9577
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8481 9537 8493 9571
rect 8527 9537 8539 9571
rect 10054 9571 10112 9577
rect 10054 9568 10066 9571
rect 8481 9531 8539 9537
rect 8864 9540 10066 9568
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 3973 9503 4031 9509
rect 3467 9472 3556 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 3528 9444 3556 9472
rect 3973 9469 3985 9503
rect 4019 9500 4031 9503
rect 4430 9500 4436 9512
rect 4019 9472 4436 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 6822 9500 6828 9512
rect 5077 9463 5135 9469
rect 5276 9472 6828 9500
rect 3510 9392 3516 9444
rect 3568 9392 3574 9444
rect 4522 9392 4528 9444
rect 4580 9392 4586 9444
rect 5092 9432 5120 9463
rect 5276 9432 5304 9472
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 5092 9404 5304 9432
rect 5629 9435 5687 9441
rect 5629 9401 5641 9435
rect 5675 9432 5687 9435
rect 7024 9432 7052 9531
rect 8205 9503 8263 9509
rect 8205 9469 8217 9503
rect 8251 9500 8263 9503
rect 8386 9500 8392 9512
rect 8251 9472 8392 9500
rect 8251 9469 8263 9472
rect 8205 9463 8263 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8496 9432 8524 9531
rect 8864 9509 8892 9540
rect 10054 9537 10066 9540
rect 10100 9537 10112 9571
rect 10054 9531 10112 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 10367 9540 10425 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 10413 9537 10425 9540
rect 10459 9568 10471 9571
rect 10686 9568 10692 9580
rect 10459 9540 10692 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 8941 9435 8999 9441
rect 8941 9432 8953 9435
rect 5675 9404 7052 9432
rect 7300 9404 8953 9432
rect 5675 9401 5687 9404
rect 5629 9395 5687 9401
rect 7300 9376 7328 9404
rect 8941 9401 8953 9404
rect 8987 9401 8999 9435
rect 8941 9395 8999 9401
rect 3050 9324 3056 9376
rect 3108 9324 3114 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3326 9364 3332 9376
rect 3191 9336 3332 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 4488 9336 6745 9364
rect 4488 9324 4494 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7282 9364 7288 9376
rect 7064 9336 7288 9364
rect 7064 9324 7070 9336
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 7524 9336 7573 9364
rect 7524 9324 7530 9336
rect 7561 9333 7573 9336
rect 7607 9333 7619 9367
rect 7561 9327 7619 9333
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 10505 9367 10563 9373
rect 10505 9364 10517 9367
rect 9088 9336 10517 9364
rect 9088 9324 9094 9336
rect 10505 9333 10517 9336
rect 10551 9333 10563 9367
rect 10505 9327 10563 9333
rect 1104 9274 10948 9296
rect 1104 9222 2180 9274
rect 2232 9222 2244 9274
rect 2296 9222 2308 9274
rect 2360 9222 2372 9274
rect 2424 9222 2436 9274
rect 2488 9222 4641 9274
rect 4693 9222 4705 9274
rect 4757 9222 4769 9274
rect 4821 9222 4833 9274
rect 4885 9222 4897 9274
rect 4949 9222 7102 9274
rect 7154 9222 7166 9274
rect 7218 9222 7230 9274
rect 7282 9222 7294 9274
rect 7346 9222 7358 9274
rect 7410 9222 9563 9274
rect 9615 9222 9627 9274
rect 9679 9222 9691 9274
rect 9743 9222 9755 9274
rect 9807 9222 9819 9274
rect 9871 9222 10948 9274
rect 1104 9200 10948 9222
rect 1946 9120 1952 9172
rect 2004 9120 2010 9172
rect 3602 9120 3608 9172
rect 3660 9120 3666 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 9214 9160 9220 9172
rect 8527 9132 9220 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 4801 9095 4859 9101
rect 4801 9061 4813 9095
rect 4847 9092 4859 9095
rect 7285 9095 7343 9101
rect 4847 9064 6316 9092
rect 4847 9061 4859 9064
rect 4801 9055 4859 9061
rect 3050 8984 3056 9036
rect 3108 8984 3114 9036
rect 4249 9027 4307 9033
rect 4249 8993 4261 9027
rect 4295 9024 4307 9027
rect 4430 9024 4436 9036
rect 4295 8996 4436 9024
rect 4295 8993 4307 8996
rect 4249 8987 4307 8993
rect 4430 8984 4436 8996
rect 4488 8984 4494 9036
rect 6288 9033 6316 9064
rect 7285 9061 7297 9095
rect 7331 9092 7343 9095
rect 7331 9064 8616 9092
rect 7331 9061 7343 9064
rect 7285 9055 7343 9061
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 8993 6331 9027
rect 6273 8987 6331 8993
rect 8113 9027 8171 9033
rect 8113 8993 8125 9027
rect 8159 9024 8171 9027
rect 8159 8996 8340 9024
rect 8159 8993 8171 8996
rect 8113 8987 8171 8993
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2222 8956 2228 8968
rect 2179 8928 2228 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 7466 8916 7472 8968
rect 7524 8916 7530 8968
rect 7558 8916 7564 8968
rect 7616 8916 7622 8968
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 4341 8891 4399 8897
rect 4341 8857 4353 8891
rect 4387 8888 4399 8891
rect 4985 8891 5043 8897
rect 4985 8888 4997 8891
rect 4387 8860 4997 8888
rect 4387 8857 4399 8860
rect 4341 8851 4399 8857
rect 4985 8857 4997 8860
rect 5031 8857 5043 8891
rect 4985 8851 5043 8857
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8888 7343 8891
rect 7650 8888 7656 8900
rect 7331 8860 7656 8888
rect 7331 8857 7343 8860
rect 7285 8851 7343 8857
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 8036 8888 8064 8919
rect 8202 8916 8208 8968
rect 8260 8916 8266 8968
rect 8312 8965 8340 8996
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 8297 8919 8355 8925
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8444 8928 8493 8956
rect 8444 8916 8450 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8588 8956 8616 9064
rect 9030 8984 9036 9036
rect 9088 8984 9094 9036
rect 9289 8959 9347 8965
rect 9289 8956 9301 8959
rect 8588 8928 9301 8956
rect 8481 8919 8539 8925
rect 9289 8925 9301 8928
rect 9335 8925 9347 8959
rect 9289 8919 9347 8925
rect 8036 8860 8340 8888
rect 8312 8832 8340 8860
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 4433 8823 4491 8829
rect 4433 8820 4445 8823
rect 3568 8792 4445 8820
rect 3568 8780 3574 8792
rect 4433 8789 4445 8792
rect 4479 8789 4491 8823
rect 4433 8783 4491 8789
rect 5718 8780 5724 8832
rect 5776 8780 5782 8832
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 10413 8823 10471 8829
rect 10413 8789 10425 8823
rect 10459 8820 10471 8823
rect 10459 8792 11008 8820
rect 10459 8789 10471 8792
rect 10413 8783 10471 8789
rect 1104 8730 10948 8752
rect 1104 8678 2840 8730
rect 2892 8678 2904 8730
rect 2956 8678 2968 8730
rect 3020 8678 3032 8730
rect 3084 8678 3096 8730
rect 3148 8678 5301 8730
rect 5353 8678 5365 8730
rect 5417 8678 5429 8730
rect 5481 8678 5493 8730
rect 5545 8678 5557 8730
rect 5609 8678 7762 8730
rect 7814 8678 7826 8730
rect 7878 8678 7890 8730
rect 7942 8678 7954 8730
rect 8006 8678 8018 8730
rect 8070 8678 10223 8730
rect 10275 8678 10287 8730
rect 10339 8678 10351 8730
rect 10403 8678 10415 8730
rect 10467 8678 10479 8730
rect 10531 8678 10948 8730
rect 1104 8656 10948 8678
rect 2222 8576 2228 8628
rect 2280 8576 2286 8628
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5626 8616 5632 8628
rect 5399 8588 5632 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5626 8576 5632 8588
rect 5684 8616 5690 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 5684 8588 5825 8616
rect 5684 8576 5690 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 10505 8619 10563 8625
rect 6227 8588 7972 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6914 8548 6920 8560
rect 5644 8520 6920 8548
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 4246 8489 4252 8492
rect 2593 8483 2651 8489
rect 2593 8449 2605 8483
rect 2639 8480 2651 8483
rect 3053 8483 3111 8489
rect 3053 8480 3065 8483
rect 2639 8452 3065 8480
rect 2639 8449 2651 8452
rect 2593 8443 2651 8449
rect 3053 8449 3065 8452
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 4240 8443 4252 8489
rect 4246 8440 4252 8443
rect 4304 8440 4310 8492
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8381 2743 8415
rect 2685 8375 2743 8381
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2700 8344 2728 8375
rect 2774 8372 2780 8424
rect 2832 8372 2838 8424
rect 3602 8372 3608 8424
rect 3660 8372 3666 8424
rect 5644 8421 5672 8520
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 7944 8557 7972 8588
rect 10505 8585 10517 8619
rect 10551 8616 10563 8619
rect 10594 8616 10600 8628
rect 10551 8588 10600 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 7377 8551 7435 8557
rect 7377 8548 7389 8551
rect 7064 8520 7389 8548
rect 7064 8508 7070 8520
rect 7377 8517 7389 8520
rect 7423 8517 7435 8551
rect 7377 8511 7435 8517
rect 7929 8551 7987 8557
rect 7929 8517 7941 8551
rect 7975 8517 7987 8551
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 7929 8511 7987 8517
rect 8036 8520 8217 8548
rect 7392 8480 7420 8511
rect 8036 8480 8064 8520
rect 8205 8517 8217 8520
rect 8251 8517 8263 8551
rect 8205 8511 8263 8517
rect 7392 8452 8064 8480
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8449 8171 8483
rect 8113 8443 8171 8449
rect 8333 8483 8391 8489
rect 8333 8449 8345 8483
rect 8379 8480 8391 8483
rect 9950 8480 9956 8492
rect 8379 8452 9956 8480
rect 8379 8449 8391 8452
rect 8333 8443 8391 8449
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 1627 8316 2728 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 3988 8276 4016 8375
rect 5718 8372 5724 8424
rect 5776 8372 5782 8424
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 7837 8415 7895 8421
rect 7616 8384 7788 8412
rect 7616 8372 7622 8384
rect 7653 8347 7711 8353
rect 7653 8313 7665 8347
rect 7699 8313 7711 8347
rect 7760 8344 7788 8384
rect 7837 8381 7849 8415
rect 7883 8412 7895 8415
rect 8128 8412 8156 8443
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 10980 8480 11008 8792
rect 10367 8452 11008 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 7883 8384 8156 8412
rect 7883 8381 7895 8384
rect 7837 8375 7895 8381
rect 7929 8347 7987 8353
rect 7929 8344 7941 8347
rect 7760 8316 7941 8344
rect 7653 8307 7711 8313
rect 7929 8313 7941 8316
rect 7975 8313 7987 8347
rect 7929 8307 7987 8313
rect 4154 8276 4160 8288
rect 3988 8248 4160 8276
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 7668 8276 7696 8307
rect 8294 8276 8300 8288
rect 7668 8248 8300 8276
rect 8294 8236 8300 8248
rect 8352 8276 8358 8288
rect 9122 8276 9128 8288
rect 8352 8248 9128 8276
rect 8352 8236 8358 8248
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 1104 8186 10948 8208
rect 1104 8134 2180 8186
rect 2232 8134 2244 8186
rect 2296 8134 2308 8186
rect 2360 8134 2372 8186
rect 2424 8134 2436 8186
rect 2488 8134 4641 8186
rect 4693 8134 4705 8186
rect 4757 8134 4769 8186
rect 4821 8134 4833 8186
rect 4885 8134 4897 8186
rect 4949 8134 7102 8186
rect 7154 8134 7166 8186
rect 7218 8134 7230 8186
rect 7282 8134 7294 8186
rect 7346 8134 7358 8186
rect 7410 8134 9563 8186
rect 9615 8134 9627 8186
rect 9679 8134 9691 8186
rect 9743 8134 9755 8186
rect 9807 8134 9819 8186
rect 9871 8134 10948 8186
rect 1104 8112 10948 8134
rect 3053 8075 3111 8081
rect 3053 8041 3065 8075
rect 3099 8072 3111 8075
rect 3602 8072 3608 8084
rect 3099 8044 3608 8072
rect 3099 8041 3111 8044
rect 3053 8035 3111 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 3973 8075 4031 8081
rect 3973 8041 3985 8075
rect 4019 8072 4031 8075
rect 4246 8072 4252 8084
rect 4019 8044 4252 8072
rect 4019 8041 4031 8044
rect 3973 8035 4031 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5629 8075 5687 8081
rect 5629 8041 5641 8075
rect 5675 8072 5687 8075
rect 5718 8072 5724 8084
rect 5675 8044 5724 8072
rect 5675 8041 5687 8044
rect 5629 8035 5687 8041
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 1670 7896 1676 7948
rect 1728 7896 1734 7948
rect 3436 7908 4384 7936
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 3436 7877 3464 7908
rect 4356 7880 4384 7908
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 4212 7840 4261 7868
rect 4212 7828 4218 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 7558 7868 7564 7880
rect 6779 7840 7564 7868
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 8110 7828 8116 7880
rect 8168 7828 8174 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 10134 7868 10140 7880
rect 9999 7840 10140 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 1946 7809 1952 7812
rect 1940 7763 1952 7809
rect 1946 7760 1952 7763
rect 2004 7760 2010 7812
rect 4494 7803 4552 7809
rect 4494 7800 4506 7803
rect 4172 7772 4506 7800
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2682 7732 2688 7744
rect 1627 7704 2688 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 4172 7732 4200 7772
rect 4494 7769 4506 7772
rect 4540 7769 4552 7803
rect 4494 7763 4552 7769
rect 3651 7704 4200 7732
rect 6549 7735 6607 7741
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 6638 7732 6644 7744
rect 6595 7704 6644 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 8665 7735 8723 7741
rect 8665 7732 8677 7735
rect 8352 7704 8677 7732
rect 8352 7692 8358 7704
rect 8665 7701 8677 7704
rect 8711 7701 8723 7735
rect 8665 7695 8723 7701
rect 10505 7735 10563 7741
rect 10505 7701 10517 7735
rect 10551 7732 10563 7735
rect 10686 7732 10692 7744
rect 10551 7704 10692 7732
rect 10551 7701 10563 7704
rect 10505 7695 10563 7701
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 1104 7642 10948 7664
rect 1104 7590 2840 7642
rect 2892 7590 2904 7642
rect 2956 7590 2968 7642
rect 3020 7590 3032 7642
rect 3084 7590 3096 7642
rect 3148 7590 5301 7642
rect 5353 7590 5365 7642
rect 5417 7590 5429 7642
rect 5481 7590 5493 7642
rect 5545 7590 5557 7642
rect 5609 7590 7762 7642
rect 7814 7590 7826 7642
rect 7878 7590 7890 7642
rect 7942 7590 7954 7642
rect 8006 7590 8018 7642
rect 8070 7590 10223 7642
rect 10275 7590 10287 7642
rect 10339 7590 10351 7642
rect 10403 7590 10415 7642
rect 10467 7590 10479 7642
rect 10531 7590 10948 7642
rect 1104 7568 10948 7590
rect 1946 7488 1952 7540
rect 2004 7488 2010 7540
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7497 2283 7531
rect 2225 7491 2283 7497
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2240 7392 2268 7491
rect 2682 7488 2688 7540
rect 2740 7488 2746 7540
rect 3786 7488 3792 7540
rect 3844 7528 3850 7540
rect 5626 7528 5632 7540
rect 3844 7500 5632 7528
rect 3844 7488 3850 7500
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 7745 7531 7803 7537
rect 7745 7497 7757 7531
rect 7791 7497 7803 7531
rect 7745 7491 7803 7497
rect 7760 7460 7788 7491
rect 8754 7488 8760 7540
rect 8812 7528 8818 7540
rect 9769 7531 9827 7537
rect 8812 7500 9628 7528
rect 8812 7488 8818 7500
rect 8110 7460 8116 7472
rect 7760 7432 8116 7460
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 9600 7460 9628 7500
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 9950 7528 9956 7540
rect 9815 7500 9956 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 9950 7488 9956 7500
rect 10008 7488 10014 7540
rect 9600 7432 9904 7460
rect 2179 7364 2268 7392
rect 2593 7395 2651 7401
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 3418 7392 3424 7404
rect 2639 7364 3424 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 6638 7401 6644 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5776 7364 5825 7392
rect 5776 7352 5782 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 6632 7392 6644 7401
rect 6599 7364 6644 7392
rect 5813 7355 5871 7361
rect 6632 7355 6644 7364
rect 6638 7352 6644 7355
rect 6696 7352 6702 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8128 7392 8156 7420
rect 7975 7364 8156 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9876 7401 9904 7432
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 2777 7327 2835 7333
rect 2777 7324 2789 7327
rect 2740 7296 2789 7324
rect 2740 7284 2746 7296
rect 2777 7293 2789 7296
rect 2823 7293 2835 7327
rect 2777 7287 2835 7293
rect 6362 7284 6368 7336
rect 6420 7284 6426 7336
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8662 7324 8668 7336
rect 8159 7296 8668 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8662 7284 8668 7296
rect 8720 7284 8726 7336
rect 8846 7284 8852 7336
rect 8904 7284 8910 7336
rect 8938 7284 8944 7336
rect 8996 7333 9002 7336
rect 8996 7327 9024 7333
rect 9012 7293 9024 7327
rect 8996 7287 9024 7293
rect 8996 7284 9002 7287
rect 8570 7216 8576 7268
rect 8628 7216 8634 7268
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 2590 7188 2596 7200
rect 1627 7160 2596 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 3881 7191 3939 7197
rect 3881 7157 3893 7191
rect 3927 7188 3939 7191
rect 4154 7188 4160 7200
rect 3927 7160 4160 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 4154 7148 4160 7160
rect 4212 7148 4218 7200
rect 5258 7148 5264 7200
rect 5316 7148 5322 7200
rect 10505 7191 10563 7197
rect 10505 7157 10517 7191
rect 10551 7188 10563 7191
rect 10594 7188 10600 7200
rect 10551 7160 10600 7188
rect 10551 7157 10563 7160
rect 10505 7151 10563 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 1104 7098 10948 7120
rect 1104 7046 2180 7098
rect 2232 7046 2244 7098
rect 2296 7046 2308 7098
rect 2360 7046 2372 7098
rect 2424 7046 2436 7098
rect 2488 7046 4641 7098
rect 4693 7046 4705 7098
rect 4757 7046 4769 7098
rect 4821 7046 4833 7098
rect 4885 7046 4897 7098
rect 4949 7046 7102 7098
rect 7154 7046 7166 7098
rect 7218 7046 7230 7098
rect 7282 7046 7294 7098
rect 7346 7046 7358 7098
rect 7410 7046 9563 7098
rect 9615 7046 9627 7098
rect 9679 7046 9691 7098
rect 9743 7046 9755 7098
rect 9807 7046 9819 7098
rect 9871 7046 10948 7098
rect 1104 7024 10948 7046
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4396 6956 5181 6984
rect 4396 6944 4402 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 5169 6947 5227 6953
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7616 6956 7849 6984
rect 7616 6944 7622 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 7837 6947 7895 6953
rect 4522 6916 4528 6928
rect 4448 6888 4528 6916
rect 3326 6808 3332 6860
rect 3384 6808 3390 6860
rect 4448 6857 4476 6888
rect 4522 6876 4528 6888
rect 4580 6916 4586 6928
rect 4580 6888 5396 6916
rect 4580 6876 4586 6888
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 5258 6848 5264 6860
rect 4663 6820 5264 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 5258 6808 5264 6820
rect 5316 6808 5322 6860
rect 5368 6848 5396 6888
rect 5368 6820 6914 6848
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 1670 6780 1676 6792
rect 1627 6752 1676 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3694 6780 3700 6792
rect 3467 6752 3700 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 1854 6721 1860 6724
rect 1848 6675 1860 6721
rect 1854 6672 1860 6675
rect 1912 6672 1918 6724
rect 2976 6684 4108 6712
rect 2976 6653 3004 6684
rect 4080 6656 4108 6684
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 3053 6647 3111 6653
rect 3053 6613 3065 6647
rect 3099 6644 3111 6647
rect 3234 6644 3240 6656
rect 3099 6616 3240 6644
rect 3099 6613 3111 6616
rect 3053 6607 3111 6613
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4709 6647 4767 6653
rect 4709 6644 4721 6647
rect 4120 6616 4721 6644
rect 4120 6604 4126 6616
rect 4709 6613 4721 6616
rect 4755 6613 4767 6647
rect 4709 6607 4767 6613
rect 5077 6647 5135 6653
rect 5077 6613 5089 6647
rect 5123 6644 5135 6647
rect 5736 6644 5764 6743
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6886 6780 6914 6820
rect 8294 6808 8300 6860
rect 8352 6808 8358 6860
rect 8389 6851 8447 6857
rect 8389 6817 8401 6851
rect 8435 6817 8447 6851
rect 8389 6811 8447 6817
rect 8404 6780 8432 6811
rect 8570 6780 8576 6792
rect 6886 6752 8576 6780
rect 8570 6740 8576 6752
rect 8628 6740 8634 6792
rect 9582 6740 9588 6792
rect 9640 6780 9646 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9640 6752 10333 6780
rect 9640 6740 9646 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10594 6740 10600 6792
rect 10652 6740 10658 6792
rect 6178 6672 6184 6724
rect 6236 6712 6242 6724
rect 8205 6715 8263 6721
rect 8205 6712 8217 6715
rect 6236 6684 8217 6712
rect 6236 6672 6242 6684
rect 8205 6681 8217 6684
rect 8251 6681 8263 6715
rect 8205 6675 8263 6681
rect 10076 6715 10134 6721
rect 10076 6681 10088 6715
rect 10122 6712 10134 6715
rect 10122 6684 10456 6712
rect 10122 6681 10134 6684
rect 10076 6675 10134 6681
rect 5123 6616 5764 6644
rect 5123 6613 5135 6616
rect 5077 6607 5135 6613
rect 6270 6604 6276 6656
rect 6328 6644 6334 6656
rect 6638 6644 6644 6656
rect 6328 6616 6644 6644
rect 6328 6604 6334 6616
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 7282 6604 7288 6656
rect 7340 6604 7346 6656
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 8662 6644 8668 6656
rect 8352 6616 8668 6644
rect 8352 6604 8358 6616
rect 8662 6604 8668 6616
rect 8720 6644 8726 6656
rect 10428 6653 10456 6684
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8720 6616 8953 6644
rect 8720 6604 8726 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 10413 6647 10471 6653
rect 10413 6613 10425 6647
rect 10459 6613 10471 6647
rect 10413 6607 10471 6613
rect 1104 6554 10948 6576
rect 1104 6502 2840 6554
rect 2892 6502 2904 6554
rect 2956 6502 2968 6554
rect 3020 6502 3032 6554
rect 3084 6502 3096 6554
rect 3148 6502 5301 6554
rect 5353 6502 5365 6554
rect 5417 6502 5429 6554
rect 5481 6502 5493 6554
rect 5545 6502 5557 6554
rect 5609 6502 7762 6554
rect 7814 6502 7826 6554
rect 7878 6502 7890 6554
rect 7942 6502 7954 6554
rect 8006 6502 8018 6554
rect 8070 6502 10223 6554
rect 10275 6502 10287 6554
rect 10339 6502 10351 6554
rect 10403 6502 10415 6554
rect 10467 6502 10479 6554
rect 10531 6502 10948 6554
rect 1104 6480 10948 6502
rect 1854 6400 1860 6452
rect 1912 6400 1918 6452
rect 2133 6443 2191 6449
rect 2133 6409 2145 6443
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 2148 6304 2176 6403
rect 2590 6400 2596 6452
rect 2648 6400 2654 6452
rect 2961 6443 3019 6449
rect 2961 6409 2973 6443
rect 3007 6440 3019 6443
rect 3418 6440 3424 6452
rect 3007 6412 3424 6440
rect 3007 6409 3019 6412
rect 2961 6403 3019 6409
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 3694 6400 3700 6452
rect 3752 6400 3758 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6270 6440 6276 6452
rect 6227 6412 6276 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6546 6400 6552 6452
rect 6604 6440 6610 6452
rect 8386 6440 8392 6452
rect 6604 6412 8392 6440
rect 6604 6400 6610 6412
rect 8386 6400 8392 6412
rect 8444 6440 8450 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 8444 6412 9689 6440
rect 8444 6400 8450 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6372 2559 6375
rect 7006 6372 7012 6384
rect 2547 6344 5488 6372
rect 2547 6341 2559 6344
rect 2501 6335 2559 6341
rect 2087 6276 2176 6304
rect 3605 6307 3663 6313
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 3605 6273 3617 6307
rect 3651 6304 3663 6307
rect 4062 6304 4068 6316
rect 3651 6276 4068 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 4689 6307 4747 6313
rect 4689 6304 4701 6307
rect 4580 6276 4701 6304
rect 4580 6264 4586 6276
rect 4689 6273 4701 6276
rect 4735 6273 4747 6307
rect 4689 6267 4747 6273
rect 2682 6196 2688 6248
rect 2740 6196 2746 6248
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4246 6236 4252 6248
rect 4019 6208 4252 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4246 6196 4252 6208
rect 4304 6196 4310 6248
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6205 4491 6239
rect 5460 6236 5488 6344
rect 6012 6344 7012 6372
rect 6012 6313 6040 6344
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 7282 6332 7288 6384
rect 7340 6372 7346 6384
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 7340 6344 7849 6372
rect 7340 6332 7346 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 7837 6335 7895 6341
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6454 6264 6460 6316
rect 6512 6264 6518 6316
rect 6638 6313 6644 6316
rect 6621 6307 6644 6313
rect 6621 6273 6633 6307
rect 6621 6267 6644 6273
rect 6638 6264 6644 6267
rect 6696 6264 6702 6316
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10686 6304 10692 6316
rect 10643 6276 10692 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 6472 6236 6500 6264
rect 5460 6208 6500 6236
rect 4433 6199 4491 6205
rect 1762 6128 1768 6180
rect 1820 6168 1826 6180
rect 4154 6168 4160 6180
rect 1820 6140 4160 6168
rect 1820 6128 1826 6140
rect 4154 6128 4160 6140
rect 4212 6168 4218 6180
rect 4448 6168 4476 6199
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 9582 6236 9588 6248
rect 9364 6208 9588 6236
rect 9364 6196 9370 6208
rect 9582 6196 9588 6208
rect 9640 6196 9646 6248
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 4212 6140 4476 6168
rect 5813 6171 5871 6177
rect 4212 6128 4218 6140
rect 5813 6137 5825 6171
rect 5859 6168 5871 6171
rect 10244 6168 10272 6199
rect 5859 6140 6408 6168
rect 5859 6137 5871 6140
rect 5813 6131 5871 6137
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6100 1639 6103
rect 4430 6100 4436 6112
rect 1627 6072 4436 6100
rect 1627 6069 1639 6072
rect 1581 6063 1639 6069
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 6380 6100 6408 6140
rect 7668 6140 10272 6168
rect 7668 6100 7696 6140
rect 6380 6072 7696 6100
rect 7745 6103 7803 6109
rect 7745 6069 7757 6103
rect 7791 6100 7803 6103
rect 8478 6100 8484 6112
rect 7791 6072 8484 6100
rect 7791 6069 7803 6072
rect 7745 6063 7803 6069
rect 8478 6060 8484 6072
rect 8536 6100 8542 6112
rect 8938 6100 8944 6112
rect 8536 6072 8944 6100
rect 8536 6060 8542 6072
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 1104 6010 10948 6032
rect 1104 5958 2180 6010
rect 2232 5958 2244 6010
rect 2296 5958 2308 6010
rect 2360 5958 2372 6010
rect 2424 5958 2436 6010
rect 2488 5958 4641 6010
rect 4693 5958 4705 6010
rect 4757 5958 4769 6010
rect 4821 5958 4833 6010
rect 4885 5958 4897 6010
rect 4949 5958 7102 6010
rect 7154 5958 7166 6010
rect 7218 5958 7230 6010
rect 7282 5958 7294 6010
rect 7346 5958 7358 6010
rect 7410 5958 9563 6010
rect 9615 5958 9627 6010
rect 9679 5958 9691 6010
rect 9743 5958 9755 6010
rect 9807 5958 9819 6010
rect 9871 5958 10948 6010
rect 1104 5936 10948 5958
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 6420 5868 6776 5896
rect 6420 5856 6426 5868
rect 3605 5831 3663 5837
rect 3605 5797 3617 5831
rect 3651 5828 3663 5831
rect 4154 5828 4160 5840
rect 3651 5800 4160 5828
rect 3651 5797 3663 5800
rect 3605 5791 3663 5797
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 3053 5763 3111 5769
rect 3053 5729 3065 5763
rect 3099 5760 3111 5763
rect 3326 5760 3332 5772
rect 3099 5732 3332 5760
rect 3099 5729 3111 5732
rect 3053 5723 3111 5729
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 4430 5720 4436 5772
rect 4488 5760 4494 5772
rect 6748 5769 6776 5868
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 7064 5868 7205 5896
rect 7064 5856 7070 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 8754 5856 8760 5908
rect 8812 5856 8818 5908
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8904 5868 8953 5896
rect 8904 5856 8910 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 8570 5828 8576 5840
rect 7852 5800 8576 5828
rect 7852 5769 7880 5800
rect 8128 5769 8156 5800
rect 8570 5788 8576 5800
rect 8628 5788 8634 5840
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 4488 5732 4905 5760
rect 4488 5720 4494 5732
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5729 5135 5763
rect 5077 5723 5135 5729
rect 6733 5763 6791 5769
rect 6733 5729 6745 5763
rect 6779 5760 6791 5763
rect 7837 5763 7895 5769
rect 6779 5732 6960 5760
rect 6779 5729 6791 5732
rect 6733 5723 6791 5729
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 3234 5652 3240 5704
rect 3292 5652 3298 5704
rect 3881 5695 3939 5701
rect 3881 5661 3893 5695
rect 3927 5692 3939 5695
rect 5092 5692 5120 5723
rect 6086 5692 6092 5704
rect 3927 5664 6092 5692
rect 3927 5661 3939 5664
rect 3881 5655 3939 5661
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 3896 5624 3924 5655
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 2740 5596 3924 5624
rect 2740 5584 2746 5596
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 4801 5627 4859 5633
rect 4304 5596 4568 5624
rect 4304 5584 4310 5596
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 1627 5528 3157 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 3145 5525 3157 5528
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 3973 5559 4031 5565
rect 3973 5556 3985 5559
rect 3384 5528 3985 5556
rect 3384 5516 3390 5528
rect 3973 5525 3985 5528
rect 4019 5525 4031 5559
rect 3973 5519 4031 5525
rect 4430 5516 4436 5568
rect 4488 5516 4494 5568
rect 4540 5556 4568 5596
rect 4801 5593 4813 5627
rect 4847 5624 4859 5627
rect 5626 5624 5632 5636
rect 4847 5596 5632 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 6466 5627 6524 5633
rect 6466 5624 6478 5627
rect 6420 5596 6478 5624
rect 6420 5584 6426 5596
rect 6466 5593 6478 5596
rect 6512 5593 6524 5627
rect 6466 5587 6524 5593
rect 6932 5624 6960 5732
rect 7837 5729 7849 5763
rect 7883 5729 7895 5763
rect 7837 5723 7895 5729
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5760 8171 5763
rect 8159 5732 8193 5760
rect 8159 5729 8171 5732
rect 8113 5723 8171 5729
rect 8294 5720 8300 5772
rect 8352 5720 8358 5772
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 9364 5664 10333 5692
rect 9364 5652 9370 5664
rect 10321 5661 10333 5664
rect 10367 5661 10379 5695
rect 10321 5655 10379 5661
rect 8294 5624 8300 5636
rect 6932 5596 8300 5624
rect 5353 5559 5411 5565
rect 5353 5556 5365 5559
rect 4540 5528 5365 5556
rect 5353 5525 5365 5528
rect 5399 5556 5411 5559
rect 6178 5556 6184 5568
rect 5399 5528 6184 5556
rect 5399 5525 5411 5528
rect 5353 5519 5411 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6932 5565 6960 5596
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 8386 5584 8392 5636
rect 8444 5584 8450 5636
rect 10076 5627 10134 5633
rect 10076 5593 10088 5627
rect 10122 5624 10134 5627
rect 10410 5624 10416 5636
rect 10122 5596 10416 5624
rect 10122 5593 10134 5596
rect 10076 5587 10134 5593
rect 10410 5584 10416 5596
rect 10468 5584 10474 5636
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5525 6975 5559
rect 6917 5519 6975 5525
rect 7558 5516 7564 5568
rect 7616 5516 7622 5568
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 1104 5466 10948 5488
rect 1104 5414 2840 5466
rect 2892 5414 2904 5466
rect 2956 5414 2968 5466
rect 3020 5414 3032 5466
rect 3084 5414 3096 5466
rect 3148 5414 5301 5466
rect 5353 5414 5365 5466
rect 5417 5414 5429 5466
rect 5481 5414 5493 5466
rect 5545 5414 5557 5466
rect 5609 5414 7762 5466
rect 7814 5414 7826 5466
rect 7878 5414 7890 5466
rect 7942 5414 7954 5466
rect 8006 5414 8018 5466
rect 8070 5414 10223 5466
rect 10275 5414 10287 5466
rect 10339 5414 10351 5466
rect 10403 5414 10415 5466
rect 10467 5414 10479 5466
rect 10531 5414 10948 5466
rect 1104 5392 10948 5414
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 2032 5287 2090 5293
rect 2032 5253 2044 5287
rect 2078 5284 2090 5287
rect 3988 5284 4016 5315
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 4709 5355 4767 5361
rect 4709 5352 4721 5355
rect 4580 5324 4721 5352
rect 4580 5312 4586 5324
rect 4709 5321 4721 5324
rect 4755 5321 4767 5355
rect 4709 5315 4767 5321
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5352 5595 5355
rect 5626 5352 5632 5364
rect 5583 5324 5632 5352
rect 5583 5321 5595 5324
rect 5537 5315 5595 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 6362 5312 6368 5364
rect 6420 5312 6426 5364
rect 8846 5312 8852 5364
rect 8904 5352 8910 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 8904 5324 9321 5352
rect 8904 5312 8910 5324
rect 9309 5321 9321 5324
rect 9355 5321 9367 5355
rect 9309 5315 9367 5321
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10134 5352 10140 5364
rect 9815 5324 10140 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 2078 5256 4016 5284
rect 2078 5253 2090 5256
rect 2032 5247 2090 5253
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4525 5219 4583 5225
rect 4525 5216 4537 5219
rect 4488 5188 4537 5216
rect 4488 5176 4494 5188
rect 4525 5185 4537 5188
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 6178 5176 6184 5228
rect 6236 5176 6242 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6730 5216 6736 5228
rect 6595 5188 6736 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 8041 5219 8099 5225
rect 8041 5185 8053 5219
rect 8087 5216 8099 5219
rect 8202 5216 8208 5228
rect 8087 5188 8208 5216
rect 8087 5185 8099 5188
rect 8041 5179 8099 5185
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 9306 5216 9312 5228
rect 8352 5188 9312 5216
rect 8352 5176 8358 5188
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 10042 5216 10048 5228
rect 9447 5188 10048 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 10042 5176 10048 5188
rect 10100 5216 10106 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 10100 5188 10241 5216
rect 10100 5176 10106 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 1762 5108 1768 5160
rect 1820 5108 1826 5160
rect 3789 5151 3847 5157
rect 3789 5117 3801 5151
rect 3835 5117 3847 5151
rect 3789 5111 3847 5117
rect 3145 5083 3203 5089
rect 3145 5049 3157 5083
rect 3191 5080 3203 5083
rect 3804 5080 3832 5111
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 9125 5151 9183 5157
rect 9125 5148 9137 5151
rect 8628 5120 9137 5148
rect 8628 5108 8634 5120
rect 9125 5117 9137 5120
rect 9171 5117 9183 5151
rect 9125 5111 9183 5117
rect 10318 5108 10324 5160
rect 10376 5108 10382 5160
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 3191 5052 3832 5080
rect 3191 5049 3203 5052
rect 3145 5043 3203 5049
rect 8662 5040 8668 5092
rect 8720 5080 8726 5092
rect 9861 5083 9919 5089
rect 9861 5080 9873 5083
rect 8720 5052 9873 5080
rect 8720 5040 8726 5052
rect 9861 5049 9873 5052
rect 9907 5049 9919 5083
rect 9861 5043 9919 5049
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 2774 5012 2780 5024
rect 1627 4984 2780 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 2774 4972 2780 4984
rect 2832 4972 2838 5024
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 3237 5015 3295 5021
rect 3237 5012 3249 5015
rect 2924 4984 3249 5012
rect 2924 4972 2930 4984
rect 3237 4981 3249 4984
rect 3283 4981 3295 5015
rect 3237 4975 3295 4981
rect 6914 4972 6920 5024
rect 6972 4972 6978 5024
rect 8846 4972 8852 5024
rect 8904 5012 8910 5024
rect 10428 5012 10456 5111
rect 8904 4984 10456 5012
rect 8904 4972 8910 4984
rect 1104 4922 10948 4944
rect 1104 4870 2180 4922
rect 2232 4870 2244 4922
rect 2296 4870 2308 4922
rect 2360 4870 2372 4922
rect 2424 4870 2436 4922
rect 2488 4870 4641 4922
rect 4693 4870 4705 4922
rect 4757 4870 4769 4922
rect 4821 4870 4833 4922
rect 4885 4870 4897 4922
rect 4949 4870 7102 4922
rect 7154 4870 7166 4922
rect 7218 4870 7230 4922
rect 7282 4870 7294 4922
rect 7346 4870 7358 4922
rect 7410 4870 9563 4922
rect 9615 4870 9627 4922
rect 9679 4870 9691 4922
rect 9743 4870 9755 4922
rect 9807 4870 9819 4922
rect 9871 4870 10948 4922
rect 1104 4848 10948 4870
rect 6730 4768 6736 4820
rect 6788 4768 6794 4820
rect 6825 4811 6883 4817
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 7558 4808 7564 4820
rect 6871 4780 7564 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 2501 4743 2559 4749
rect 2501 4709 2513 4743
rect 2547 4709 2559 4743
rect 2501 4703 2559 4709
rect 5077 4743 5135 4749
rect 5077 4709 5089 4743
rect 5123 4740 5135 4743
rect 5718 4740 5724 4752
rect 5123 4712 5724 4740
rect 5123 4709 5135 4712
rect 5077 4703 5135 4709
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2516 4604 2544 4703
rect 5718 4700 5724 4712
rect 5776 4700 5782 4752
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2832 4644 2973 4672
rect 2832 4632 2838 4644
rect 2961 4641 2973 4644
rect 3007 4641 3019 4675
rect 2961 4635 3019 4641
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 3326 4672 3332 4684
rect 3191 4644 3332 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 6086 4632 6092 4684
rect 6144 4632 6150 4684
rect 2363 4576 2544 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2866 4564 2872 4616
rect 2924 4564 2930 4616
rect 4338 4564 4344 4616
rect 4396 4564 4402 4616
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5626 4604 5632 4616
rect 4939 4576 5632 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 5810 4564 5816 4616
rect 5868 4564 5874 4616
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 6840 4604 6868 4771
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7708 4780 7757 4808
rect 7708 4768 7714 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 8260 4780 8493 4808
rect 8260 4768 8266 4780
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 9306 4808 9312 4820
rect 8481 4771 8539 4777
rect 8956 4780 9312 4808
rect 6914 4632 6920 4684
rect 6972 4672 6978 4684
rect 7377 4675 7435 4681
rect 7377 4672 7389 4675
rect 6972 4644 7389 4672
rect 6972 4632 6978 4644
rect 7377 4641 7389 4644
rect 7423 4641 7435 4675
rect 7377 4635 7435 4641
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 8478 4672 8484 4684
rect 8435 4644 8484 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8478 4632 8484 4644
rect 8536 4632 8542 4684
rect 8956 4681 8984 4780
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 10318 4768 10324 4820
rect 10376 4808 10382 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 10376 4780 10425 4808
rect 10376 4768 10382 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 10413 4771 10471 4777
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4641 8999 4675
rect 8941 4635 8999 4641
rect 6411 4576 6868 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 8662 4564 8668 4616
rect 8720 4564 8726 4616
rect 10594 4564 10600 4616
rect 10652 4564 10658 4616
rect 9208 4539 9266 4545
rect 9208 4505 9220 4539
rect 9254 4536 9266 4539
rect 9582 4536 9588 4548
rect 9254 4508 9588 4536
rect 9254 4505 9266 4508
rect 9208 4499 9266 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 2130 4428 2136 4480
rect 2188 4428 2194 4480
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 3789 4471 3847 4477
rect 3789 4468 3801 4471
rect 3292 4440 3801 4468
rect 3292 4428 3298 4440
rect 3789 4437 3801 4440
rect 3835 4437 3847 4471
rect 3789 4431 3847 4437
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4468 4859 4471
rect 5074 4468 5080 4480
rect 4847 4440 5080 4468
rect 4847 4437 4859 4440
rect 4801 4431 4859 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5166 4428 5172 4480
rect 5224 4428 5230 4480
rect 6270 4428 6276 4480
rect 6328 4428 6334 4480
rect 10134 4428 10140 4480
rect 10192 4468 10198 4480
rect 10321 4471 10379 4477
rect 10321 4468 10333 4471
rect 10192 4440 10333 4468
rect 10192 4428 10198 4440
rect 10321 4437 10333 4440
rect 10367 4437 10379 4471
rect 10321 4431 10379 4437
rect 1104 4378 10948 4400
rect 1104 4326 2840 4378
rect 2892 4326 2904 4378
rect 2956 4326 2968 4378
rect 3020 4326 3032 4378
rect 3084 4326 3096 4378
rect 3148 4326 5301 4378
rect 5353 4326 5365 4378
rect 5417 4326 5429 4378
rect 5481 4326 5493 4378
rect 5545 4326 5557 4378
rect 5609 4326 7762 4378
rect 7814 4326 7826 4378
rect 7878 4326 7890 4378
rect 7942 4326 7954 4378
rect 8006 4326 8018 4378
rect 8070 4326 10223 4378
rect 10275 4326 10287 4378
rect 10339 4326 10351 4378
rect 10403 4326 10415 4378
rect 10467 4326 10479 4378
rect 10531 4326 10948 4378
rect 1104 4304 10948 4326
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 4709 4267 4767 4273
rect 4709 4264 4721 4267
rect 4672 4236 4721 4264
rect 4672 4224 4678 4236
rect 4709 4233 4721 4236
rect 4755 4233 4767 4267
rect 4709 4227 4767 4233
rect 5077 4267 5135 4273
rect 5077 4233 5089 4267
rect 5123 4264 5135 4267
rect 5166 4264 5172 4276
rect 5123 4236 5172 4264
rect 5123 4233 5135 4236
rect 5077 4227 5135 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 6365 4267 6423 4273
rect 6365 4264 6377 4267
rect 5684 4236 6377 4264
rect 5684 4224 5690 4236
rect 6365 4233 6377 4236
rect 6411 4233 6423 4267
rect 6365 4227 6423 4233
rect 9582 4224 9588 4276
rect 9640 4224 9646 4276
rect 9861 4267 9919 4273
rect 9861 4233 9873 4267
rect 9907 4264 9919 4267
rect 10042 4264 10048 4276
rect 9907 4236 10048 4264
rect 9907 4233 9919 4236
rect 9861 4227 9919 4233
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 2032 4199 2090 4205
rect 2032 4165 2044 4199
rect 2078 4196 2090 4199
rect 2130 4196 2136 4208
rect 2078 4168 2136 4196
rect 2078 4165 2090 4168
rect 2032 4159 2090 4165
rect 2130 4156 2136 4168
rect 2188 4156 2194 4208
rect 9125 4199 9183 4205
rect 9125 4165 9137 4199
rect 9171 4196 9183 4199
rect 9950 4196 9956 4208
rect 9171 4168 9956 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 9950 4156 9956 4168
rect 10008 4156 10014 4208
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3602 4128 3608 4140
rect 3559 4100 3608 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 6227 4100 6745 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4128 8355 4131
rect 8938 4128 8944 4140
rect 8343 4100 8944 4128
rect 8343 4097 8355 4100
rect 8297 4091 8355 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 9508 4100 9781 4128
rect 1762 4020 1768 4072
rect 1820 4020 1826 4072
rect 3786 4020 3792 4072
rect 3844 4020 3850 4072
rect 5166 4020 5172 4072
rect 5224 4020 5230 4072
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4029 5411 4063
rect 5353 4023 5411 4029
rect 3145 3995 3203 4001
rect 3145 3961 3157 3995
rect 3191 3992 3203 3995
rect 4338 3992 4344 4004
rect 3191 3964 4344 3992
rect 3191 3961 3203 3964
rect 3145 3955 3203 3961
rect 4338 3952 4344 3964
rect 4396 3952 4402 4004
rect 5368 3992 5396 4023
rect 5626 4020 5632 4072
rect 5684 4020 5690 4072
rect 6086 4020 6092 4072
rect 6144 4060 6150 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6144 4032 6837 4060
rect 6144 4020 6150 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4029 7067 4063
rect 7009 4023 7067 4029
rect 6914 3992 6920 4004
rect 5368 3964 6920 3992
rect 6914 3952 6920 3964
rect 6972 3992 6978 4004
rect 7024 3992 7052 4023
rect 7558 4020 7564 4072
rect 7616 4060 7622 4072
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7616 4032 7757 4060
rect 7616 4020 7622 4032
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4060 8263 4063
rect 8478 4060 8484 4072
rect 8251 4032 8484 4060
rect 8251 4029 8263 4032
rect 8205 4023 8263 4029
rect 8128 3992 8156 4023
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8846 4020 8852 4072
rect 8904 4020 8910 4072
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 8864 3992 8892 4020
rect 6972 3964 8892 3992
rect 6972 3952 6978 3964
rect 3694 3884 3700 3936
rect 3752 3884 3758 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 4433 3927 4491 3933
rect 4433 3924 4445 3927
rect 4028 3896 4445 3924
rect 4028 3884 4034 3896
rect 4433 3893 4445 3896
rect 4479 3893 4491 3927
rect 4433 3887 4491 3893
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7193 3927 7251 3933
rect 7193 3924 7205 3927
rect 7064 3896 7205 3924
rect 7064 3884 7070 3896
rect 7193 3893 7205 3896
rect 7239 3893 7251 3927
rect 7193 3887 7251 3893
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 8628 3896 8677 3924
rect 8628 3884 8634 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 9048 3924 9076 4023
rect 9508 4001 9536 4100
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 10192 4100 10425 4128
rect 10192 4088 10198 4100
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 9493 3995 9551 4001
rect 9493 3961 9505 3995
rect 9539 3961 9551 3995
rect 9493 3955 9551 3961
rect 10410 3924 10416 3936
rect 9048 3896 10416 3924
rect 8665 3887 8723 3893
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 1104 3834 10948 3856
rect 1104 3782 2180 3834
rect 2232 3782 2244 3834
rect 2296 3782 2308 3834
rect 2360 3782 2372 3834
rect 2424 3782 2436 3834
rect 2488 3782 4641 3834
rect 4693 3782 4705 3834
rect 4757 3782 4769 3834
rect 4821 3782 4833 3834
rect 4885 3782 4897 3834
rect 4949 3782 7102 3834
rect 7154 3782 7166 3834
rect 7218 3782 7230 3834
rect 7282 3782 7294 3834
rect 7346 3782 7358 3834
rect 7410 3782 9563 3834
rect 9615 3782 9627 3834
rect 9679 3782 9691 3834
rect 9743 3782 9755 3834
rect 9807 3782 9819 3834
rect 9871 3782 10948 3834
rect 1104 3760 10948 3782
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 3786 3720 3792 3732
rect 3651 3692 3792 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5810 3720 5816 3732
rect 5215 3692 5816 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 6825 3723 6883 3729
rect 6825 3689 6837 3723
rect 6871 3720 6883 3723
rect 7558 3720 7564 3732
rect 6871 3692 7564 3720
rect 6871 3689 6883 3692
rect 6825 3683 6883 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8938 3680 8944 3732
rect 8996 3680 9002 3732
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9950 3720 9956 3732
rect 9723 3692 9956 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10410 3680 10416 3732
rect 10468 3680 10474 3732
rect 8297 3655 8355 3661
rect 8297 3621 8309 3655
rect 8343 3652 8355 3655
rect 8343 3624 9536 3652
rect 8343 3621 8355 3624
rect 8297 3615 8355 3621
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 9508 3593 9536 3624
rect 9493 3587 9551 3593
rect 1820 3556 2268 3584
rect 1820 3544 1826 3556
rect 1946 3476 1952 3528
rect 2004 3476 2010 3528
rect 2240 3525 2268 3556
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 2271 3488 3801 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 3789 3485 3801 3488
rect 3835 3516 3847 3519
rect 4798 3516 4804 3528
rect 3835 3488 4804 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5445 3519 5503 3525
rect 5445 3485 5457 3519
rect 5491 3516 5503 3519
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 5491 3488 6929 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 6917 3485 6929 3488
rect 6963 3516 6975 3519
rect 8294 3516 8300 3528
rect 6963 3488 8300 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9640 3488 10241 3516
rect 9640 3476 9646 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10229 3479 10287 3485
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 2470 3451 2528 3457
rect 2470 3448 2482 3451
rect 2148 3420 2482 3448
rect 2148 3389 2176 3420
rect 2470 3417 2482 3420
rect 2516 3417 2528 3451
rect 2470 3411 2528 3417
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 5718 3457 5724 3460
rect 4034 3451 4092 3457
rect 4034 3448 4046 3451
rect 3752 3420 4046 3448
rect 3752 3408 3758 3420
rect 4034 3417 4046 3420
rect 4080 3417 4092 3451
rect 5712 3448 5724 3457
rect 5679 3420 5724 3448
rect 4034 3411 4092 3417
rect 5712 3411 5724 3420
rect 5718 3408 5724 3411
rect 5776 3408 5782 3460
rect 7184 3451 7242 3457
rect 7184 3417 7196 3451
rect 7230 3448 7242 3451
rect 7650 3448 7656 3460
rect 7230 3420 7656 3448
rect 7230 3417 7242 3420
rect 7184 3411 7242 3417
rect 7650 3408 7656 3420
rect 7708 3408 7714 3460
rect 2133 3383 2191 3389
rect 2133 3349 2145 3383
rect 2179 3349 2191 3383
rect 2133 3343 2191 3349
rect 8386 3340 8392 3392
rect 8444 3340 8450 3392
rect 1104 3290 10948 3312
rect 1104 3238 2840 3290
rect 2892 3238 2904 3290
rect 2956 3238 2968 3290
rect 3020 3238 3032 3290
rect 3084 3238 3096 3290
rect 3148 3238 5301 3290
rect 5353 3238 5365 3290
rect 5417 3238 5429 3290
rect 5481 3238 5493 3290
rect 5545 3238 5557 3290
rect 5609 3238 7762 3290
rect 7814 3238 7826 3290
rect 7878 3238 7890 3290
rect 7942 3238 7954 3290
rect 8006 3238 8018 3290
rect 8070 3238 10223 3290
rect 10275 3238 10287 3290
rect 10339 3238 10351 3290
rect 10403 3238 10415 3290
rect 10467 3238 10479 3290
rect 10531 3238 10948 3290
rect 1104 3216 10948 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2004 3148 2697 3176
rect 2004 3136 2010 3148
rect 2685 3145 2697 3148
rect 2731 3145 2743 3179
rect 2685 3139 2743 3145
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3234 3176 3240 3188
rect 3099 3148 3240 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 3602 3136 3608 3188
rect 3660 3136 3666 3188
rect 3970 3136 3976 3188
rect 4028 3136 4034 3188
rect 5626 3136 5632 3188
rect 5684 3176 5690 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5684 3148 6193 3176
rect 5684 3136 5690 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 7006 3136 7012 3188
rect 7064 3176 7070 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 7064 3148 7205 3176
rect 7064 3136 7070 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 7561 3179 7619 3185
rect 7561 3145 7573 3179
rect 7607 3145 7619 3179
rect 7561 3139 7619 3145
rect 4065 3111 4123 3117
rect 4065 3077 4077 3111
rect 4111 3108 4123 3111
rect 4154 3108 4160 3120
rect 4111 3080 4160 3108
rect 4111 3077 4123 3080
rect 4065 3071 4123 3077
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 5074 3117 5080 3120
rect 5068 3108 5080 3117
rect 5035 3080 5080 3108
rect 5068 3071 5080 3080
rect 5074 3068 5080 3071
rect 5132 3068 5138 3120
rect 4798 3000 4804 3052
rect 4856 3000 4862 3052
rect 6914 3040 6920 3052
rect 4908 3012 6920 3040
rect 3142 2932 3148 2984
rect 3200 2932 3206 2984
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 3384 2944 4261 2972
rect 3384 2932 3390 2944
rect 4249 2941 4261 2944
rect 4295 2972 4307 2975
rect 4908 2972 4936 3012
rect 6914 3000 6920 3012
rect 6972 3040 6978 3052
rect 7576 3040 7604 3139
rect 7650 3136 7656 3188
rect 7708 3136 7714 3188
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 9401 3179 9459 3185
rect 9401 3145 9413 3179
rect 9447 3176 9459 3179
rect 9582 3176 9588 3188
rect 9447 3148 9588 3176
rect 9447 3145 9459 3148
rect 9401 3139 9459 3145
rect 9582 3136 9588 3148
rect 9640 3136 9646 3188
rect 8312 3108 8340 3136
rect 8036 3080 8340 3108
rect 8036 3049 8064 3080
rect 8386 3068 8392 3120
rect 8444 3068 8450 3120
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 6972 3012 7052 3040
rect 7576 3012 7849 3040
rect 6972 3000 6978 3012
rect 7024 2981 7052 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 8021 3043 8079 3049
rect 8021 3009 8033 3043
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 8288 3043 8346 3049
rect 8288 3009 8300 3043
rect 8334 3040 8346 3043
rect 8404 3040 8432 3068
rect 8334 3012 8432 3040
rect 8334 3009 8346 3012
rect 8288 3003 8346 3009
rect 4295 2944 4936 2972
rect 7009 2975 7067 2981
rect 4295 2941 4307 2944
rect 4249 2935 4307 2941
rect 7009 2941 7021 2975
rect 7055 2941 7067 2975
rect 7009 2935 7067 2941
rect 7098 2932 7104 2984
rect 7156 2932 7162 2984
rect 1104 2746 10948 2768
rect 1104 2694 2180 2746
rect 2232 2694 2244 2746
rect 2296 2694 2308 2746
rect 2360 2694 2372 2746
rect 2424 2694 2436 2746
rect 2488 2694 4641 2746
rect 4693 2694 4705 2746
rect 4757 2694 4769 2746
rect 4821 2694 4833 2746
rect 4885 2694 4897 2746
rect 4949 2694 7102 2746
rect 7154 2694 7166 2746
rect 7218 2694 7230 2746
rect 7282 2694 7294 2746
rect 7346 2694 7358 2746
rect 7410 2694 9563 2746
rect 9615 2694 9627 2746
rect 9679 2694 9691 2746
rect 9743 2694 9755 2746
rect 9807 2694 9819 2746
rect 9871 2694 10948 2746
rect 1104 2672 10948 2694
rect 3142 2592 3148 2644
rect 3200 2632 3206 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 3200 2604 3341 2632
rect 3200 2592 3206 2604
rect 3329 2601 3341 2604
rect 3375 2601 3387 2635
rect 3329 2595 3387 2601
rect 4154 2592 4160 2644
rect 4212 2592 4218 2644
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 5224 2604 5273 2632
rect 5224 2592 5230 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 6086 2592 6092 2644
rect 6144 2592 6150 2644
rect 6270 2592 6276 2644
rect 6328 2632 6334 2644
rect 6549 2635 6607 2641
rect 6549 2632 6561 2635
rect 6328 2604 6561 2632
rect 6328 2592 6334 2604
rect 6549 2601 6561 2604
rect 6595 2601 6607 2635
rect 6549 2595 6607 2601
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7193 2635 7251 2641
rect 7193 2632 7205 2635
rect 7064 2604 7205 2632
rect 7064 2592 7070 2604
rect 7193 2601 7205 2604
rect 7239 2601 7251 2635
rect 7193 2595 7251 2601
rect 8478 2592 8484 2644
rect 8536 2592 8542 2644
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 3292 2400 3525 2428
rect 3292 2388 3298 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5224 2400 5457 2428
rect 5224 2388 5230 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5868 2400 5917 2428
rect 5868 2388 5874 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6512 2400 6745 2428
rect 6512 2388 6518 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7156 2400 7389 2428
rect 7156 2388 7162 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 8444 2400 8677 2428
rect 8444 2388 8450 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 1104 2202 10948 2224
rect 1104 2150 2840 2202
rect 2892 2150 2904 2202
rect 2956 2150 2968 2202
rect 3020 2150 3032 2202
rect 3084 2150 3096 2202
rect 3148 2150 5301 2202
rect 5353 2150 5365 2202
rect 5417 2150 5429 2202
rect 5481 2150 5493 2202
rect 5545 2150 5557 2202
rect 5609 2150 7762 2202
rect 7814 2150 7826 2202
rect 7878 2150 7890 2202
rect 7942 2150 7954 2202
rect 8006 2150 8018 2202
rect 8070 2150 10223 2202
rect 10275 2150 10287 2202
rect 10339 2150 10351 2202
rect 10403 2150 10415 2202
rect 10467 2150 10479 2202
rect 10531 2150 10948 2202
rect 1104 2128 10948 2150
<< via1 >>
rect 2840 11942 2892 11994
rect 2904 11942 2956 11994
rect 2968 11942 3020 11994
rect 3032 11942 3084 11994
rect 3096 11942 3148 11994
rect 5301 11942 5353 11994
rect 5365 11942 5417 11994
rect 5429 11942 5481 11994
rect 5493 11942 5545 11994
rect 5557 11942 5609 11994
rect 7762 11942 7814 11994
rect 7826 11942 7878 11994
rect 7890 11942 7942 11994
rect 7954 11942 8006 11994
rect 8018 11942 8070 11994
rect 10223 11942 10275 11994
rect 10287 11942 10339 11994
rect 10351 11942 10403 11994
rect 10415 11942 10467 11994
rect 10479 11942 10531 11994
rect 5172 11704 5224 11756
rect 4528 11636 4580 11688
rect 7656 11704 7708 11756
rect 4160 11568 4212 11620
rect 4344 11500 4396 11552
rect 7564 11500 7616 11552
rect 2180 11398 2232 11450
rect 2244 11398 2296 11450
rect 2308 11398 2360 11450
rect 2372 11398 2424 11450
rect 2436 11398 2488 11450
rect 4641 11398 4693 11450
rect 4705 11398 4757 11450
rect 4769 11398 4821 11450
rect 4833 11398 4885 11450
rect 4897 11398 4949 11450
rect 7102 11398 7154 11450
rect 7166 11398 7218 11450
rect 7230 11398 7282 11450
rect 7294 11398 7346 11450
rect 7358 11398 7410 11450
rect 9563 11398 9615 11450
rect 9627 11398 9679 11450
rect 9691 11398 9743 11450
rect 9755 11398 9807 11450
rect 9819 11398 9871 11450
rect 5172 11296 5224 11348
rect 4436 11160 4488 11212
rect 2504 11092 2556 11144
rect 3332 11092 3384 11144
rect 4252 11092 4304 11144
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 7564 11092 7616 11144
rect 7656 11092 7708 11144
rect 4896 11024 4948 11076
rect 6184 11024 6236 11076
rect 2228 10999 2280 11008
rect 2228 10965 2237 10999
rect 2237 10965 2271 10999
rect 2271 10965 2280 10999
rect 2228 10956 2280 10965
rect 6276 10999 6328 11008
rect 6276 10965 6285 10999
rect 6285 10965 6319 10999
rect 6319 10965 6328 10999
rect 6276 10956 6328 10965
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 8944 11024 8996 11076
rect 8208 10956 8260 11008
rect 2840 10854 2892 10906
rect 2904 10854 2956 10906
rect 2968 10854 3020 10906
rect 3032 10854 3084 10906
rect 3096 10854 3148 10906
rect 5301 10854 5353 10906
rect 5365 10854 5417 10906
rect 5429 10854 5481 10906
rect 5493 10854 5545 10906
rect 5557 10854 5609 10906
rect 7762 10854 7814 10906
rect 7826 10854 7878 10906
rect 7890 10854 7942 10906
rect 7954 10854 8006 10906
rect 8018 10854 8070 10906
rect 10223 10854 10275 10906
rect 10287 10854 10339 10906
rect 10351 10854 10403 10906
rect 10415 10854 10467 10906
rect 10479 10854 10531 10906
rect 3332 10795 3384 10804
rect 3332 10761 3341 10795
rect 3341 10761 3375 10795
rect 3375 10761 3384 10795
rect 3332 10752 3384 10761
rect 5172 10752 5224 10804
rect 6092 10752 6144 10804
rect 7656 10752 7708 10804
rect 848 10616 900 10668
rect 1676 10616 1728 10668
rect 2228 10659 2280 10668
rect 2228 10625 2262 10659
rect 2262 10625 2280 10659
rect 2228 10616 2280 10625
rect 4160 10684 4212 10736
rect 4896 10684 4948 10736
rect 6184 10727 6236 10736
rect 6184 10693 6193 10727
rect 6193 10693 6227 10727
rect 6227 10693 6236 10727
rect 6184 10684 6236 10693
rect 6276 10684 6328 10736
rect 8944 10727 8996 10736
rect 8944 10693 8962 10727
rect 8962 10693 8996 10727
rect 8944 10684 8996 10693
rect 6460 10616 6512 10668
rect 3608 10591 3660 10600
rect 3608 10557 3617 10591
rect 3617 10557 3651 10591
rect 3651 10557 3660 10591
rect 3608 10548 3660 10557
rect 5172 10548 5224 10600
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 10416 10548 10468 10600
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 7012 10412 7064 10464
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 7840 10412 7892 10421
rect 2180 10310 2232 10362
rect 2244 10310 2296 10362
rect 2308 10310 2360 10362
rect 2372 10310 2424 10362
rect 2436 10310 2488 10362
rect 4641 10310 4693 10362
rect 4705 10310 4757 10362
rect 4769 10310 4821 10362
rect 4833 10310 4885 10362
rect 4897 10310 4949 10362
rect 7102 10310 7154 10362
rect 7166 10310 7218 10362
rect 7230 10310 7282 10362
rect 7294 10310 7346 10362
rect 7358 10310 7410 10362
rect 9563 10310 9615 10362
rect 9627 10310 9679 10362
rect 9691 10310 9743 10362
rect 9755 10310 9807 10362
rect 9819 10310 9871 10362
rect 2504 10208 2556 10260
rect 5172 10251 5224 10260
rect 5172 10217 5181 10251
rect 5181 10217 5215 10251
rect 5215 10217 5224 10251
rect 5172 10208 5224 10217
rect 1584 10072 1636 10124
rect 2688 10004 2740 10056
rect 3608 10072 3660 10124
rect 4344 10004 4396 10056
rect 7012 10004 7064 10056
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 3608 9868 3660 9920
rect 6368 9936 6420 9988
rect 6184 9868 6236 9920
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 10416 10251 10468 10260
rect 10416 10217 10425 10251
rect 10425 10217 10459 10251
rect 10459 10217 10468 10251
rect 10416 10208 10468 10217
rect 7748 10140 7800 10192
rect 7656 10072 7708 10124
rect 8576 10140 8628 10192
rect 10692 10072 10744 10124
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7840 9936 7892 9988
rect 8576 9936 8628 9988
rect 9220 9936 9272 9988
rect 8300 9868 8352 9920
rect 2840 9766 2892 9818
rect 2904 9766 2956 9818
rect 2968 9766 3020 9818
rect 3032 9766 3084 9818
rect 3096 9766 3148 9818
rect 5301 9766 5353 9818
rect 5365 9766 5417 9818
rect 5429 9766 5481 9818
rect 5493 9766 5545 9818
rect 5557 9766 5609 9818
rect 7762 9766 7814 9818
rect 7826 9766 7878 9818
rect 7890 9766 7942 9818
rect 7954 9766 8006 9818
rect 8018 9766 8070 9818
rect 10223 9766 10275 9818
rect 10287 9766 10339 9818
rect 10351 9766 10403 9818
rect 10415 9766 10467 9818
rect 10479 9766 10531 9818
rect 5172 9664 5224 9716
rect 4252 9596 4304 9648
rect 5080 9596 5132 9648
rect 8300 9664 8352 9716
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 1952 9571 2004 9580
rect 1952 9537 1986 9571
rect 1986 9537 2004 9571
rect 1952 9528 2004 9537
rect 3332 9528 3384 9580
rect 3608 9528 3660 9580
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 8208 9596 8260 9648
rect 4436 9460 4488 9512
rect 3516 9392 3568 9444
rect 4528 9435 4580 9444
rect 4528 9401 4537 9435
rect 4537 9401 4571 9435
rect 4571 9401 4580 9435
rect 4528 9392 4580 9401
rect 6828 9460 6880 9512
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 10692 9528 10744 9580
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 3332 9324 3384 9376
rect 4436 9324 4488 9376
rect 7012 9324 7064 9376
rect 7288 9367 7340 9376
rect 7288 9333 7297 9367
rect 7297 9333 7331 9367
rect 7331 9333 7340 9367
rect 7288 9324 7340 9333
rect 7472 9324 7524 9376
rect 9036 9324 9088 9376
rect 2180 9222 2232 9274
rect 2244 9222 2296 9274
rect 2308 9222 2360 9274
rect 2372 9222 2424 9274
rect 2436 9222 2488 9274
rect 4641 9222 4693 9274
rect 4705 9222 4757 9274
rect 4769 9222 4821 9274
rect 4833 9222 4885 9274
rect 4897 9222 4949 9274
rect 7102 9222 7154 9274
rect 7166 9222 7218 9274
rect 7230 9222 7282 9274
rect 7294 9222 7346 9274
rect 7358 9222 7410 9274
rect 9563 9222 9615 9274
rect 9627 9222 9679 9274
rect 9691 9222 9743 9274
rect 9755 9222 9807 9274
rect 9819 9222 9871 9274
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 9220 9120 9272 9172
rect 3056 9027 3108 9036
rect 3056 8993 3065 9027
rect 3065 8993 3099 9027
rect 3099 8993 3108 9027
rect 3056 8984 3108 8993
rect 4436 8984 4488 9036
rect 2228 8916 2280 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 7564 8959 7616 8968
rect 7564 8925 7573 8959
rect 7573 8925 7607 8959
rect 7607 8925 7616 8959
rect 7564 8916 7616 8925
rect 7656 8848 7708 8900
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8392 8916 8444 8968
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 3516 8780 3568 8832
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 8300 8780 8352 8832
rect 2840 8678 2892 8730
rect 2904 8678 2956 8730
rect 2968 8678 3020 8730
rect 3032 8678 3084 8730
rect 3096 8678 3148 8730
rect 5301 8678 5353 8730
rect 5365 8678 5417 8730
rect 5429 8678 5481 8730
rect 5493 8678 5545 8730
rect 5557 8678 5609 8730
rect 7762 8678 7814 8730
rect 7826 8678 7878 8730
rect 7890 8678 7942 8730
rect 7954 8678 8006 8730
rect 8018 8678 8070 8730
rect 10223 8678 10275 8730
rect 10287 8678 10339 8730
rect 10351 8678 10403 8730
rect 10415 8678 10467 8730
rect 10479 8678 10531 8730
rect 2228 8619 2280 8628
rect 2228 8585 2237 8619
rect 2237 8585 2271 8619
rect 2271 8585 2280 8619
rect 2228 8576 2280 8585
rect 5632 8576 5684 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 4252 8483 4304 8492
rect 4252 8449 4286 8483
rect 4286 8449 4304 8483
rect 4252 8440 4304 8449
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 6920 8508 6972 8560
rect 7012 8508 7064 8560
rect 10600 8576 10652 8628
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 7564 8372 7616 8424
rect 9956 8440 10008 8492
rect 4160 8236 4212 8288
rect 8300 8236 8352 8288
rect 9128 8236 9180 8288
rect 2180 8134 2232 8186
rect 2244 8134 2296 8186
rect 2308 8134 2360 8186
rect 2372 8134 2424 8186
rect 2436 8134 2488 8186
rect 4641 8134 4693 8186
rect 4705 8134 4757 8186
rect 4769 8134 4821 8186
rect 4833 8134 4885 8186
rect 4897 8134 4949 8186
rect 7102 8134 7154 8186
rect 7166 8134 7218 8186
rect 7230 8134 7282 8186
rect 7294 8134 7346 8186
rect 7358 8134 7410 8186
rect 9563 8134 9615 8186
rect 9627 8134 9679 8186
rect 9691 8134 9743 8186
rect 9755 8134 9807 8186
rect 9819 8134 9871 8186
rect 3608 8032 3660 8084
rect 4252 8032 4304 8084
rect 5724 8032 5776 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 848 7828 900 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4160 7828 4212 7880
rect 4344 7828 4396 7880
rect 7564 7828 7616 7880
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 10140 7828 10192 7880
rect 1952 7803 2004 7812
rect 1952 7769 1986 7803
rect 1986 7769 2004 7803
rect 1952 7760 2004 7769
rect 2688 7692 2740 7744
rect 6644 7692 6696 7744
rect 8300 7692 8352 7744
rect 10692 7692 10744 7744
rect 2840 7590 2892 7642
rect 2904 7590 2956 7642
rect 2968 7590 3020 7642
rect 3032 7590 3084 7642
rect 3096 7590 3148 7642
rect 5301 7590 5353 7642
rect 5365 7590 5417 7642
rect 5429 7590 5481 7642
rect 5493 7590 5545 7642
rect 5557 7590 5609 7642
rect 7762 7590 7814 7642
rect 7826 7590 7878 7642
rect 7890 7590 7942 7642
rect 7954 7590 8006 7642
rect 8018 7590 8070 7642
rect 10223 7590 10275 7642
rect 10287 7590 10339 7642
rect 10351 7590 10403 7642
rect 10415 7590 10467 7642
rect 10479 7590 10531 7642
rect 1952 7531 2004 7540
rect 1952 7497 1961 7531
rect 1961 7497 1995 7531
rect 1995 7497 2004 7531
rect 1952 7488 2004 7497
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2688 7531 2740 7540
rect 2688 7497 2697 7531
rect 2697 7497 2731 7531
rect 2731 7497 2740 7531
rect 2688 7488 2740 7497
rect 3792 7488 3844 7540
rect 5632 7488 5684 7540
rect 8760 7488 8812 7540
rect 8116 7420 8168 7472
rect 9956 7488 10008 7540
rect 3424 7352 3476 7404
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5724 7352 5776 7404
rect 6644 7395 6696 7404
rect 6644 7361 6678 7395
rect 6678 7361 6696 7395
rect 6644 7352 6696 7361
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 2688 7284 2740 7336
rect 6368 7327 6420 7336
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 8668 7284 8720 7336
rect 8852 7327 8904 7336
rect 8852 7293 8861 7327
rect 8861 7293 8895 7327
rect 8895 7293 8904 7327
rect 8852 7284 8904 7293
rect 8944 7327 8996 7336
rect 8944 7293 8978 7327
rect 8978 7293 8996 7327
rect 8944 7284 8996 7293
rect 8576 7259 8628 7268
rect 8576 7225 8585 7259
rect 8585 7225 8619 7259
rect 8619 7225 8628 7259
rect 8576 7216 8628 7225
rect 2596 7148 2648 7200
rect 4160 7148 4212 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 10600 7148 10652 7200
rect 2180 7046 2232 7098
rect 2244 7046 2296 7098
rect 2308 7046 2360 7098
rect 2372 7046 2424 7098
rect 2436 7046 2488 7098
rect 4641 7046 4693 7098
rect 4705 7046 4757 7098
rect 4769 7046 4821 7098
rect 4833 7046 4885 7098
rect 4897 7046 4949 7098
rect 7102 7046 7154 7098
rect 7166 7046 7218 7098
rect 7230 7046 7282 7098
rect 7294 7046 7346 7098
rect 7358 7046 7410 7098
rect 9563 7046 9615 7098
rect 9627 7046 9679 7098
rect 9691 7046 9743 7098
rect 9755 7046 9807 7098
rect 9819 7046 9871 7098
rect 4344 6944 4396 6996
rect 7564 6944 7616 6996
rect 3332 6851 3384 6860
rect 3332 6817 3341 6851
rect 3341 6817 3375 6851
rect 3375 6817 3384 6851
rect 3332 6808 3384 6817
rect 4528 6876 4580 6928
rect 5264 6808 5316 6860
rect 1676 6740 1728 6792
rect 3700 6740 3752 6792
rect 1860 6715 1912 6724
rect 1860 6681 1894 6715
rect 1894 6681 1912 6715
rect 1860 6672 1912 6681
rect 3240 6604 3292 6656
rect 4068 6604 4120 6656
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 8300 6851 8352 6860
rect 8300 6817 8309 6851
rect 8309 6817 8343 6851
rect 8343 6817 8352 6851
rect 8300 6808 8352 6817
rect 8576 6740 8628 6792
rect 9588 6740 9640 6792
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 6184 6672 6236 6724
rect 6276 6604 6328 6656
rect 6644 6604 6696 6656
rect 7288 6647 7340 6656
rect 7288 6613 7297 6647
rect 7297 6613 7331 6647
rect 7331 6613 7340 6647
rect 7288 6604 7340 6613
rect 8300 6604 8352 6656
rect 8668 6604 8720 6656
rect 2840 6502 2892 6554
rect 2904 6502 2956 6554
rect 2968 6502 3020 6554
rect 3032 6502 3084 6554
rect 3096 6502 3148 6554
rect 5301 6502 5353 6554
rect 5365 6502 5417 6554
rect 5429 6502 5481 6554
rect 5493 6502 5545 6554
rect 5557 6502 5609 6554
rect 7762 6502 7814 6554
rect 7826 6502 7878 6554
rect 7890 6502 7942 6554
rect 7954 6502 8006 6554
rect 8018 6502 8070 6554
rect 10223 6502 10275 6554
rect 10287 6502 10339 6554
rect 10351 6502 10403 6554
rect 10415 6502 10467 6554
rect 10479 6502 10531 6554
rect 1860 6443 1912 6452
rect 1860 6409 1869 6443
rect 1869 6409 1903 6443
rect 1903 6409 1912 6443
rect 1860 6400 1912 6409
rect 848 6264 900 6316
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 3424 6400 3476 6452
rect 3700 6443 3752 6452
rect 3700 6409 3709 6443
rect 3709 6409 3743 6443
rect 3743 6409 3752 6443
rect 3700 6400 3752 6409
rect 6276 6400 6328 6452
rect 6552 6400 6604 6452
rect 8392 6400 8444 6452
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4528 6264 4580 6316
rect 2688 6239 2740 6248
rect 2688 6205 2697 6239
rect 2697 6205 2731 6239
rect 2731 6205 2740 6239
rect 2688 6196 2740 6205
rect 4252 6196 4304 6248
rect 7012 6332 7064 6384
rect 7288 6332 7340 6384
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6460 6264 6512 6316
rect 6644 6307 6696 6316
rect 6644 6273 6667 6307
rect 6667 6273 6696 6307
rect 6644 6264 6696 6273
rect 10692 6264 10744 6316
rect 1768 6128 1820 6180
rect 4160 6128 4212 6180
rect 9312 6196 9364 6248
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 4436 6060 4488 6112
rect 8484 6060 8536 6112
rect 8944 6060 8996 6112
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 2180 5958 2232 6010
rect 2244 5958 2296 6010
rect 2308 5958 2360 6010
rect 2372 5958 2424 6010
rect 2436 5958 2488 6010
rect 4641 5958 4693 6010
rect 4705 5958 4757 6010
rect 4769 5958 4821 6010
rect 4833 5958 4885 6010
rect 4897 5958 4949 6010
rect 7102 5958 7154 6010
rect 7166 5958 7218 6010
rect 7230 5958 7282 6010
rect 7294 5958 7346 6010
rect 7358 5958 7410 6010
rect 9563 5958 9615 6010
rect 9627 5958 9679 6010
rect 9691 5958 9743 6010
rect 9755 5958 9807 6010
rect 9819 5958 9871 6010
rect 6368 5856 6420 5908
rect 4160 5788 4212 5840
rect 3332 5720 3384 5772
rect 4436 5720 4488 5772
rect 7012 5856 7064 5908
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 8852 5856 8904 5908
rect 8576 5788 8628 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 2688 5584 2740 5636
rect 6092 5652 6144 5704
rect 4252 5584 4304 5636
rect 3332 5516 3384 5568
rect 4436 5559 4488 5568
rect 4436 5525 4445 5559
rect 4445 5525 4479 5559
rect 4479 5525 4488 5559
rect 4436 5516 4488 5525
rect 5632 5584 5684 5636
rect 6368 5584 6420 5636
rect 8300 5763 8352 5772
rect 8300 5729 8309 5763
rect 8309 5729 8343 5763
rect 8343 5729 8352 5763
rect 8300 5720 8352 5729
rect 9312 5652 9364 5704
rect 6184 5516 6236 5568
rect 8300 5584 8352 5636
rect 8392 5627 8444 5636
rect 8392 5593 8401 5627
rect 8401 5593 8435 5627
rect 8435 5593 8444 5627
rect 8392 5584 8444 5593
rect 10416 5584 10468 5636
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 2840 5414 2892 5466
rect 2904 5414 2956 5466
rect 2968 5414 3020 5466
rect 3032 5414 3084 5466
rect 3096 5414 3148 5466
rect 5301 5414 5353 5466
rect 5365 5414 5417 5466
rect 5429 5414 5481 5466
rect 5493 5414 5545 5466
rect 5557 5414 5609 5466
rect 7762 5414 7814 5466
rect 7826 5414 7878 5466
rect 7890 5414 7942 5466
rect 7954 5414 8006 5466
rect 8018 5414 8070 5466
rect 10223 5414 10275 5466
rect 10287 5414 10339 5466
rect 10351 5414 10403 5466
rect 10415 5414 10467 5466
rect 10479 5414 10531 5466
rect 4528 5312 4580 5364
rect 5632 5312 5684 5364
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 8852 5312 8904 5364
rect 10140 5312 10192 5364
rect 848 5176 900 5228
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 4436 5176 4488 5228
rect 6184 5219 6236 5228
rect 6184 5185 6193 5219
rect 6193 5185 6227 5219
rect 6227 5185 6236 5219
rect 6184 5176 6236 5185
rect 6736 5176 6788 5228
rect 8208 5176 8260 5228
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 9312 5176 9364 5228
rect 10048 5176 10100 5228
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 8576 5108 8628 5160
rect 10324 5151 10376 5160
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 8668 5040 8720 5092
rect 2780 4972 2832 5024
rect 2872 4972 2924 5024
rect 6920 5015 6972 5024
rect 6920 4981 6929 5015
rect 6929 4981 6963 5015
rect 6963 4981 6972 5015
rect 6920 4972 6972 4981
rect 8852 4972 8904 5024
rect 2180 4870 2232 4922
rect 2244 4870 2296 4922
rect 2308 4870 2360 4922
rect 2372 4870 2424 4922
rect 2436 4870 2488 4922
rect 4641 4870 4693 4922
rect 4705 4870 4757 4922
rect 4769 4870 4821 4922
rect 4833 4870 4885 4922
rect 4897 4870 4949 4922
rect 7102 4870 7154 4922
rect 7166 4870 7218 4922
rect 7230 4870 7282 4922
rect 7294 4870 7346 4922
rect 7358 4870 7410 4922
rect 9563 4870 9615 4922
rect 9627 4870 9679 4922
rect 9691 4870 9743 4922
rect 9755 4870 9807 4922
rect 9819 4870 9871 4922
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 5724 4700 5776 4752
rect 2780 4632 2832 4684
rect 3332 4632 3384 4684
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 4344 4607 4396 4616
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 5632 4564 5684 4616
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 7564 4768 7616 4820
rect 7656 4768 7708 4820
rect 8208 4768 8260 4820
rect 6920 4632 6972 4684
rect 8484 4632 8536 4684
rect 9312 4768 9364 4820
rect 10324 4768 10376 4820
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10643 4607
rect 10643 4573 10652 4607
rect 10600 4564 10652 4573
rect 9588 4496 9640 4548
rect 2136 4471 2188 4480
rect 2136 4437 2145 4471
rect 2145 4437 2179 4471
rect 2179 4437 2188 4471
rect 2136 4428 2188 4437
rect 3240 4428 3292 4480
rect 5080 4428 5132 4480
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 6276 4471 6328 4480
rect 6276 4437 6285 4471
rect 6285 4437 6319 4471
rect 6319 4437 6328 4471
rect 6276 4428 6328 4437
rect 10140 4428 10192 4480
rect 2840 4326 2892 4378
rect 2904 4326 2956 4378
rect 2968 4326 3020 4378
rect 3032 4326 3084 4378
rect 3096 4326 3148 4378
rect 5301 4326 5353 4378
rect 5365 4326 5417 4378
rect 5429 4326 5481 4378
rect 5493 4326 5545 4378
rect 5557 4326 5609 4378
rect 7762 4326 7814 4378
rect 7826 4326 7878 4378
rect 7890 4326 7942 4378
rect 7954 4326 8006 4378
rect 8018 4326 8070 4378
rect 10223 4326 10275 4378
rect 10287 4326 10339 4378
rect 10351 4326 10403 4378
rect 10415 4326 10467 4378
rect 10479 4326 10531 4378
rect 4620 4224 4672 4276
rect 5172 4224 5224 4276
rect 5632 4224 5684 4276
rect 9588 4267 9640 4276
rect 9588 4233 9597 4267
rect 9597 4233 9631 4267
rect 9631 4233 9640 4267
rect 9588 4224 9640 4233
rect 10048 4224 10100 4276
rect 2136 4156 2188 4208
rect 9956 4156 10008 4208
rect 3608 4088 3660 4140
rect 8944 4088 8996 4140
rect 1768 4063 1820 4072
rect 1768 4029 1777 4063
rect 1777 4029 1811 4063
rect 1811 4029 1820 4063
rect 1768 4020 1820 4029
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 5172 4020 5224 4029
rect 4344 3952 4396 4004
rect 5632 4063 5684 4072
rect 5632 4029 5641 4063
rect 5641 4029 5675 4063
rect 5675 4029 5684 4063
rect 5632 4020 5684 4029
rect 6092 4020 6144 4072
rect 6920 3952 6972 4004
rect 7564 4020 7616 4072
rect 8484 4020 8536 4072
rect 8852 4063 8904 4072
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 3976 3884 4028 3936
rect 7012 3884 7064 3936
rect 8576 3884 8628 3936
rect 10140 4088 10192 4140
rect 10416 3884 10468 3936
rect 2180 3782 2232 3834
rect 2244 3782 2296 3834
rect 2308 3782 2360 3834
rect 2372 3782 2424 3834
rect 2436 3782 2488 3834
rect 4641 3782 4693 3834
rect 4705 3782 4757 3834
rect 4769 3782 4821 3834
rect 4833 3782 4885 3834
rect 4897 3782 4949 3834
rect 7102 3782 7154 3834
rect 7166 3782 7218 3834
rect 7230 3782 7282 3834
rect 7294 3782 7346 3834
rect 7358 3782 7410 3834
rect 9563 3782 9615 3834
rect 9627 3782 9679 3834
rect 9691 3782 9743 3834
rect 9755 3782 9807 3834
rect 9819 3782 9871 3834
rect 3792 3680 3844 3732
rect 5816 3680 5868 3732
rect 7564 3680 7616 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 9956 3680 10008 3732
rect 10416 3723 10468 3732
rect 10416 3689 10425 3723
rect 10425 3689 10459 3723
rect 10459 3689 10468 3723
rect 10416 3680 10468 3689
rect 1768 3544 1820 3596
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 4804 3476 4856 3528
rect 8300 3476 8352 3528
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 9588 3476 9640 3528
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 3700 3408 3752 3460
rect 5724 3451 5776 3460
rect 5724 3417 5758 3451
rect 5758 3417 5776 3451
rect 5724 3408 5776 3417
rect 7656 3408 7708 3460
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 2840 3238 2892 3290
rect 2904 3238 2956 3290
rect 2968 3238 3020 3290
rect 3032 3238 3084 3290
rect 3096 3238 3148 3290
rect 5301 3238 5353 3290
rect 5365 3238 5417 3290
rect 5429 3238 5481 3290
rect 5493 3238 5545 3290
rect 5557 3238 5609 3290
rect 7762 3238 7814 3290
rect 7826 3238 7878 3290
rect 7890 3238 7942 3290
rect 7954 3238 8006 3290
rect 8018 3238 8070 3290
rect 10223 3238 10275 3290
rect 10287 3238 10339 3290
rect 10351 3238 10403 3290
rect 10415 3238 10467 3290
rect 10479 3238 10531 3290
rect 1952 3136 2004 3188
rect 3240 3136 3292 3188
rect 3608 3179 3660 3188
rect 3608 3145 3617 3179
rect 3617 3145 3651 3179
rect 3651 3145 3660 3179
rect 3608 3136 3660 3145
rect 3976 3179 4028 3188
rect 3976 3145 3985 3179
rect 3985 3145 4019 3179
rect 4019 3145 4028 3179
rect 3976 3136 4028 3145
rect 5632 3136 5684 3188
rect 7012 3136 7064 3188
rect 4160 3068 4212 3120
rect 5080 3111 5132 3120
rect 5080 3077 5114 3111
rect 5114 3077 5132 3111
rect 5080 3068 5132 3077
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 3148 2975 3200 2984
rect 3148 2941 3157 2975
rect 3157 2941 3191 2975
rect 3191 2941 3200 2975
rect 3148 2932 3200 2941
rect 3332 2975 3384 2984
rect 3332 2941 3341 2975
rect 3341 2941 3375 2975
rect 3375 2941 3384 2975
rect 3332 2932 3384 2941
rect 6920 3000 6972 3052
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 8300 3136 8352 3188
rect 9588 3136 9640 3188
rect 8392 3068 8444 3120
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 2180 2694 2232 2746
rect 2244 2694 2296 2746
rect 2308 2694 2360 2746
rect 2372 2694 2424 2746
rect 2436 2694 2488 2746
rect 4641 2694 4693 2746
rect 4705 2694 4757 2746
rect 4769 2694 4821 2746
rect 4833 2694 4885 2746
rect 4897 2694 4949 2746
rect 7102 2694 7154 2746
rect 7166 2694 7218 2746
rect 7230 2694 7282 2746
rect 7294 2694 7346 2746
rect 7358 2694 7410 2746
rect 9563 2694 9615 2746
rect 9627 2694 9679 2746
rect 9691 2694 9743 2746
rect 9755 2694 9807 2746
rect 9819 2694 9871 2746
rect 3148 2592 3200 2644
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 5172 2592 5224 2644
rect 6092 2635 6144 2644
rect 6092 2601 6101 2635
rect 6101 2601 6135 2635
rect 6135 2601 6144 2635
rect 6092 2592 6144 2601
rect 6276 2592 6328 2644
rect 7012 2592 7064 2644
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 3240 2388 3292 2440
rect 3884 2388 3936 2440
rect 5172 2388 5224 2440
rect 5816 2388 5868 2440
rect 6460 2388 6512 2440
rect 7104 2388 7156 2440
rect 8392 2388 8444 2440
rect 2840 2150 2892 2202
rect 2904 2150 2956 2202
rect 2968 2150 3020 2202
rect 3032 2150 3084 2202
rect 3096 2150 3148 2202
rect 5301 2150 5353 2202
rect 5365 2150 5417 2202
rect 5429 2150 5481 2202
rect 5493 2150 5545 2202
rect 5557 2150 5609 2202
rect 7762 2150 7814 2202
rect 7826 2150 7878 2202
rect 7890 2150 7942 2202
rect 7954 2150 8006 2202
rect 8018 2150 8070 2202
rect 10223 2150 10275 2202
rect 10287 2150 10339 2202
rect 10351 2150 10403 2202
rect 10415 2150 10467 2202
rect 10479 2150 10531 2202
<< metal2 >>
rect 7746 13466 7802 14266
rect 7760 12186 7788 13466
rect 7668 12158 7788 12186
rect 2840 11996 3148 12005
rect 2840 11994 2846 11996
rect 2902 11994 2926 11996
rect 2982 11994 3006 11996
rect 3062 11994 3086 11996
rect 3142 11994 3148 11996
rect 2902 11942 2904 11994
rect 3084 11942 3086 11994
rect 2840 11940 2846 11942
rect 2902 11940 2926 11942
rect 2982 11940 3006 11942
rect 3062 11940 3086 11942
rect 3142 11940 3148 11942
rect 2840 11931 3148 11940
rect 5301 11996 5609 12005
rect 5301 11994 5307 11996
rect 5363 11994 5387 11996
rect 5443 11994 5467 11996
rect 5523 11994 5547 11996
rect 5603 11994 5609 11996
rect 5363 11942 5365 11994
rect 5545 11942 5547 11994
rect 5301 11940 5307 11942
rect 5363 11940 5387 11942
rect 5443 11940 5467 11942
rect 5523 11940 5547 11942
rect 5603 11940 5609 11942
rect 5301 11931 5609 11940
rect 7668 11762 7696 12158
rect 7762 11996 8070 12005
rect 7762 11994 7768 11996
rect 7824 11994 7848 11996
rect 7904 11994 7928 11996
rect 7984 11994 8008 11996
rect 8064 11994 8070 11996
rect 7824 11942 7826 11994
rect 8006 11942 8008 11994
rect 7762 11940 7768 11942
rect 7824 11940 7848 11942
rect 7904 11940 7928 11942
rect 7984 11940 8008 11942
rect 8064 11940 8070 11942
rect 7762 11931 8070 11940
rect 10223 11996 10531 12005
rect 10223 11994 10229 11996
rect 10285 11994 10309 11996
rect 10365 11994 10389 11996
rect 10445 11994 10469 11996
rect 10525 11994 10531 11996
rect 10285 11942 10287 11994
rect 10467 11942 10469 11994
rect 10223 11940 10229 11942
rect 10285 11940 10309 11942
rect 10365 11940 10389 11942
rect 10445 11940 10469 11942
rect 10525 11940 10531 11942
rect 10223 11931 10531 11940
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4160 11620 4212 11626
rect 4160 11562 4212 11568
rect 2180 11452 2488 11461
rect 2180 11450 2186 11452
rect 2242 11450 2266 11452
rect 2322 11450 2346 11452
rect 2402 11450 2426 11452
rect 2482 11450 2488 11452
rect 2242 11398 2244 11450
rect 2424 11398 2426 11450
rect 2180 11396 2186 11398
rect 2242 11396 2266 11398
rect 2322 11396 2346 11398
rect 2402 11396 2426 11398
rect 2482 11396 2488 11398
rect 2180 11387 2488 11396
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2240 10674 2268 10950
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 860 10441 888 10610
rect 1584 10464 1636 10470
rect 846 10432 902 10441
rect 1584 10406 1636 10412
rect 846 10367 902 10376
rect 1596 10130 1624 10406
rect 1584 10124 1636 10130
rect 1584 10066 1636 10072
rect 1688 9586 1716 10610
rect 2180 10364 2488 10373
rect 2180 10362 2186 10364
rect 2242 10362 2266 10364
rect 2322 10362 2346 10364
rect 2402 10362 2426 10364
rect 2482 10362 2488 10364
rect 2242 10310 2244 10362
rect 2424 10310 2426 10362
rect 2180 10308 2186 10310
rect 2242 10308 2266 10310
rect 2322 10308 2346 10310
rect 2402 10308 2426 10310
rect 2482 10308 2488 10310
rect 2180 10299 2488 10308
rect 2516 10266 2544 11086
rect 2840 10908 3148 10917
rect 2840 10906 2846 10908
rect 2902 10906 2926 10908
rect 2982 10906 3006 10908
rect 3062 10906 3086 10908
rect 3142 10906 3148 10908
rect 2902 10854 2904 10906
rect 3084 10854 3086 10906
rect 2840 10852 2846 10854
rect 2902 10852 2926 10854
rect 2982 10852 3006 10854
rect 3062 10852 3086 10854
rect 3142 10852 3148 10854
rect 2840 10843 3148 10852
rect 3344 10810 3372 11086
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1688 7954 1716 9522
rect 1964 9178 1992 9522
rect 2180 9276 2488 9285
rect 2180 9274 2186 9276
rect 2242 9274 2266 9276
rect 2322 9274 2346 9276
rect 2402 9274 2426 9276
rect 2482 9274 2488 9276
rect 2242 9222 2244 9274
rect 2424 9222 2426 9274
rect 2180 9220 2186 9222
rect 2242 9220 2266 9222
rect 2322 9220 2346 9222
rect 2402 9220 2426 9222
rect 2482 9220 2488 9222
rect 2180 9211 2488 9220
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2240 8634 2268 8910
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2700 8378 2728 9998
rect 2840 9820 3148 9829
rect 2840 9818 2846 9820
rect 2902 9818 2926 9820
rect 2982 9818 3006 9820
rect 3062 9818 3086 9820
rect 3142 9818 3148 9820
rect 2902 9766 2904 9818
rect 3084 9766 3086 9818
rect 2840 9764 2846 9766
rect 2902 9764 2926 9766
rect 2982 9764 3006 9766
rect 3062 9764 3086 9766
rect 3142 9764 3148 9766
rect 2840 9755 3148 9764
rect 3344 9586 3372 10746
rect 4172 10742 4200 11562
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3620 10130 3648 10542
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9586 3648 9862
rect 4264 9654 4292 11086
rect 4356 10062 4384 11494
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3068 9042 3096 9318
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2840 8732 3148 8741
rect 2840 8730 2846 8732
rect 2902 8730 2926 8732
rect 2982 8730 3006 8732
rect 3062 8730 3086 8732
rect 3142 8730 3148 8732
rect 2902 8678 2904 8730
rect 3084 8678 3086 8730
rect 2840 8676 2846 8678
rect 2902 8676 2926 8678
rect 2982 8676 3006 8678
rect 3062 8676 3086 8678
rect 3142 8676 3148 8678
rect 2840 8667 3148 8676
rect 2780 8424 2832 8430
rect 2608 8372 2780 8378
rect 2608 8366 2832 8372
rect 2608 8350 2820 8366
rect 2180 8188 2488 8197
rect 2180 8186 2186 8188
rect 2242 8186 2266 8188
rect 2322 8186 2346 8188
rect 2402 8186 2426 8188
rect 2482 8186 2488 8188
rect 2242 8134 2244 8186
rect 2424 8134 2426 8186
rect 2180 8132 2186 8134
rect 2242 8132 2266 8134
rect 2322 8132 2346 8134
rect 2402 8132 2426 8134
rect 2482 8132 2488 8134
rect 2180 8123 2488 8132
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6905 1440 7346
rect 1688 6914 1716 7890
rect 1952 7812 2004 7818
rect 1952 7754 2004 7760
rect 1964 7546 1992 7754
rect 1952 7540 2004 7546
rect 1952 7482 2004 7488
rect 2608 7426 2636 8350
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2700 7546 2728 7686
rect 2840 7644 3148 7653
rect 2840 7642 2846 7644
rect 2902 7642 2926 7644
rect 2982 7642 3006 7644
rect 3062 7642 3086 7644
rect 3142 7642 3148 7644
rect 2902 7590 2904 7642
rect 3084 7590 3086 7642
rect 2840 7588 2846 7590
rect 2902 7588 2926 7590
rect 2982 7588 3006 7590
rect 3062 7588 3086 7590
rect 3142 7588 3148 7590
rect 2840 7579 3148 7588
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2608 7398 2728 7426
rect 2700 7342 2728 7398
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2180 7100 2488 7109
rect 2180 7098 2186 7100
rect 2242 7098 2266 7100
rect 2322 7098 2346 7100
rect 2402 7098 2426 7100
rect 2482 7098 2488 7100
rect 2242 7046 2244 7098
rect 2424 7046 2426 7098
rect 2180 7044 2186 7046
rect 2242 7044 2266 7046
rect 2322 7044 2346 7046
rect 2402 7044 2426 7046
rect 2482 7044 2488 7046
rect 2180 7035 2488 7044
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 1688 6886 1808 6914
rect 1688 6798 1716 6886
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1780 6186 1808 6886
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6458 1900 6666
rect 2608 6458 2636 7142
rect 1860 6452 1912 6458
rect 1860 6394 1912 6400
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2700 6254 2728 7278
rect 3344 6866 3372 9318
rect 3528 8838 3556 9386
rect 3620 9178 3648 9522
rect 4448 9518 4476 11154
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4448 9382 4476 9454
rect 4540 9450 4568 11630
rect 4641 11452 4949 11461
rect 4641 11450 4647 11452
rect 4703 11450 4727 11452
rect 4783 11450 4807 11452
rect 4863 11450 4887 11452
rect 4943 11450 4949 11452
rect 4703 11398 4705 11450
rect 4885 11398 4887 11450
rect 4641 11396 4647 11398
rect 4703 11396 4727 11398
rect 4783 11396 4807 11398
rect 4863 11396 4887 11398
rect 4943 11396 4949 11398
rect 4641 11387 4949 11396
rect 5184 11354 5212 11698
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7102 11452 7410 11461
rect 7102 11450 7108 11452
rect 7164 11450 7188 11452
rect 7244 11450 7268 11452
rect 7324 11450 7348 11452
rect 7404 11450 7410 11452
rect 7164 11398 7166 11450
rect 7346 11398 7348 11450
rect 7102 11396 7108 11398
rect 7164 11396 7188 11398
rect 7244 11396 7268 11398
rect 7324 11396 7348 11398
rect 7404 11396 7410 11398
rect 7102 11387 7410 11396
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 7576 11150 7604 11494
rect 9563 11452 9871 11461
rect 9563 11450 9569 11452
rect 9625 11450 9649 11452
rect 9705 11450 9729 11452
rect 9785 11450 9809 11452
rect 9865 11450 9871 11452
rect 9625 11398 9627 11450
rect 9807 11398 9809 11450
rect 9563 11396 9569 11398
rect 9625 11396 9649 11398
rect 9705 11396 9729 11398
rect 9785 11396 9809 11398
rect 9865 11396 9871 11398
rect 9563 11387 9871 11396
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4908 10742 4936 11018
rect 5184 10810 5212 11086
rect 5301 10908 5609 10917
rect 5301 10906 5307 10908
rect 5363 10906 5387 10908
rect 5443 10906 5467 10908
rect 5523 10906 5547 10908
rect 5603 10906 5609 10908
rect 5363 10854 5365 10906
rect 5545 10854 5547 10906
rect 5301 10852 5307 10854
rect 5363 10852 5387 10854
rect 5443 10852 5467 10854
rect 5523 10852 5547 10854
rect 5603 10852 5609 10854
rect 5301 10843 5609 10852
rect 6104 10810 6132 11086
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 4896 10736 4948 10742
rect 5184 10690 5212 10746
rect 6196 10742 6224 11018
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6288 10742 6316 10950
rect 4896 10678 4948 10684
rect 5092 10662 5212 10690
rect 6184 10736 6236 10742
rect 6184 10678 6236 10684
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 4641 10364 4949 10373
rect 4641 10362 4647 10364
rect 4703 10362 4727 10364
rect 4783 10362 4807 10364
rect 4863 10362 4887 10364
rect 4943 10362 4949 10364
rect 4703 10310 4705 10362
rect 4885 10310 4887 10362
rect 4641 10308 4647 10310
rect 4703 10308 4727 10310
rect 4783 10308 4807 10310
rect 4863 10308 4887 10310
rect 4943 10308 4949 10310
rect 4641 10299 4949 10308
rect 5092 9654 5120 10662
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10266 5212 10542
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5184 9722 5212 10202
rect 6196 9926 6224 10678
rect 6472 10674 6500 11086
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6380 9994 6408 10542
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10062 7052 10406
rect 7102 10364 7410 10373
rect 7102 10362 7108 10364
rect 7164 10362 7188 10364
rect 7244 10362 7268 10364
rect 7324 10362 7348 10364
rect 7404 10362 7410 10364
rect 7164 10310 7166 10362
rect 7346 10310 7348 10362
rect 7102 10308 7108 10310
rect 7164 10308 7188 10310
rect 7244 10308 7268 10310
rect 7324 10308 7348 10310
rect 7404 10308 7410 10310
rect 7102 10299 7410 10308
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7576 10010 7604 11086
rect 7668 10810 7696 11086
rect 7762 10908 8070 10917
rect 7762 10906 7768 10908
rect 7824 10906 7848 10908
rect 7904 10906 7928 10908
rect 7984 10906 8008 10908
rect 8064 10906 8070 10908
rect 7824 10854 7826 10906
rect 8006 10854 8008 10906
rect 7762 10852 7768 10854
rect 7824 10852 7848 10854
rect 7904 10852 7928 10854
rect 7984 10852 8008 10854
rect 8064 10852 8070 10854
rect 7762 10843 8070 10852
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7668 10130 7696 10746
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7760 10010 7788 10134
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 5301 9820 5609 9829
rect 5301 9818 5307 9820
rect 5363 9818 5387 9820
rect 5443 9818 5467 9820
rect 5523 9818 5547 9820
rect 5603 9818 5609 9820
rect 5363 9766 5365 9818
rect 5545 9766 5547 9818
rect 5301 9764 5307 9766
rect 5363 9764 5387 9766
rect 5443 9764 5467 9766
rect 5523 9764 5547 9766
rect 5603 9764 5609 9766
rect 5301 9755 5609 9764
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 4448 9042 4476 9318
rect 4641 9276 4949 9285
rect 4641 9274 4647 9276
rect 4703 9274 4727 9276
rect 4783 9274 4807 9276
rect 4863 9274 4887 9276
rect 4943 9274 4949 9276
rect 4703 9222 4705 9274
rect 4885 9222 4887 9274
rect 4641 9220 4647 9222
rect 4703 9220 4727 9222
rect 4783 9220 4807 9222
rect 4863 9220 4887 9222
rect 4943 9220 4949 9222
rect 4641 9211 4949 9220
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8650 3556 8774
rect 3528 8622 3648 8650
rect 3620 8430 3648 8622
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3620 8090 3648 8366
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 4172 7886 4200 8230
rect 4264 8090 4292 8434
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 3804 7546 3832 7822
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 2840 6556 3148 6565
rect 2840 6554 2846 6556
rect 2902 6554 2926 6556
rect 2982 6554 3006 6556
rect 3062 6554 3086 6556
rect 3142 6554 3148 6556
rect 2902 6502 2904 6554
rect 3084 6502 3086 6554
rect 2840 6500 2846 6502
rect 2902 6500 2926 6502
rect 2982 6500 3006 6502
rect 3062 6500 3086 6502
rect 3142 6500 3148 6502
rect 2840 6491 3148 6500
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 1780 5166 1808 6122
rect 2180 6012 2488 6021
rect 2180 6010 2186 6012
rect 2242 6010 2266 6012
rect 2322 6010 2346 6012
rect 2402 6010 2426 6012
rect 2482 6010 2488 6012
rect 2242 5958 2244 6010
rect 2424 5958 2426 6010
rect 2180 5956 2186 5958
rect 2242 5956 2266 5958
rect 2322 5956 2346 5958
rect 2402 5956 2426 5958
rect 2482 5956 2488 5958
rect 2180 5947 2488 5956
rect 2700 5642 2728 6190
rect 3252 5710 3280 6598
rect 3436 6458 3464 7346
rect 4172 7206 4200 7822
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3712 6458 3740 6734
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 4080 6322 4108 6598
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4172 6186 4200 7142
rect 4356 7002 4384 7822
rect 4448 7018 4476 8978
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5301 8732 5609 8741
rect 5301 8730 5307 8732
rect 5363 8730 5387 8732
rect 5443 8730 5467 8732
rect 5523 8730 5547 8732
rect 5603 8730 5609 8732
rect 5363 8678 5365 8730
rect 5545 8678 5547 8730
rect 5301 8676 5307 8678
rect 5363 8676 5387 8678
rect 5443 8676 5467 8678
rect 5523 8676 5547 8678
rect 5603 8676 5609 8678
rect 5301 8667 5609 8676
rect 5644 8634 5672 8910
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5736 8514 5764 8774
rect 5644 8486 5764 8514
rect 4641 8188 4949 8197
rect 4641 8186 4647 8188
rect 4703 8186 4727 8188
rect 4783 8186 4807 8188
rect 4863 8186 4887 8188
rect 4943 8186 4949 8188
rect 4703 8134 4705 8186
rect 4885 8134 4887 8186
rect 4641 8132 4647 8134
rect 4703 8132 4727 8134
rect 4783 8132 4807 8134
rect 4863 8132 4887 8134
rect 4943 8132 4949 8134
rect 4641 8123 4949 8132
rect 5301 7644 5609 7653
rect 5301 7642 5307 7644
rect 5363 7642 5387 7644
rect 5443 7642 5467 7644
rect 5523 7642 5547 7644
rect 5603 7642 5609 7644
rect 5363 7590 5365 7642
rect 5545 7590 5547 7642
rect 5301 7588 5307 7590
rect 5363 7588 5387 7590
rect 5443 7588 5467 7590
rect 5523 7588 5547 7590
rect 5603 7588 5609 7590
rect 5301 7579 5609 7588
rect 5644 7546 5672 8486
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8090 5764 8366
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5736 7410 5764 8026
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 4641 7100 4949 7109
rect 4641 7098 4647 7100
rect 4703 7098 4727 7100
rect 4783 7098 4807 7100
rect 4863 7098 4887 7100
rect 4943 7098 4949 7100
rect 4703 7046 4705 7098
rect 4885 7046 4887 7098
rect 4641 7044 4647 7046
rect 4703 7044 4727 7046
rect 4783 7044 4807 7046
rect 4863 7044 4887 7046
rect 4943 7044 4949 7046
rect 4641 7035 4949 7044
rect 5184 7041 5212 7346
rect 6380 7342 6408 9930
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9586 6960 9862
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 9512 6880 9518
rect 7024 9466 7052 9998
rect 6880 9460 7052 9466
rect 6828 9454 7052 9460
rect 6840 9438 7052 9454
rect 6932 8566 6960 9438
rect 7300 9382 7328 9998
rect 7576 9982 7788 10010
rect 7852 9994 7880 10406
rect 8128 10266 8156 11086
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8220 10266 8248 10950
rect 8956 10742 8984 11018
rect 10223 10908 10531 10917
rect 10223 10906 10229 10908
rect 10285 10906 10309 10908
rect 10365 10906 10389 10908
rect 10445 10906 10469 10908
rect 10525 10906 10531 10908
rect 10285 10854 10287 10906
rect 10467 10854 10469 10906
rect 10223 10852 10229 10854
rect 10285 10852 10309 10854
rect 10365 10852 10389 10854
rect 10445 10852 10469 10854
rect 10525 10852 10531 10854
rect 10223 10843 10531 10852
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 9563 10364 9871 10373
rect 9563 10362 9569 10364
rect 9625 10362 9649 10364
rect 9705 10362 9729 10364
rect 9785 10362 9809 10364
rect 9865 10362 9871 10364
rect 9625 10310 9627 10362
rect 9807 10310 9809 10362
rect 9563 10308 9569 10310
rect 9625 10308 9649 10310
rect 9705 10308 9729 10310
rect 9785 10308 9809 10310
rect 9865 10308 9871 10310
rect 9563 10299 9871 10308
rect 10428 10266 10456 10542
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 7840 9988 7892 9994
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7024 8566 7052 9318
rect 7102 9276 7410 9285
rect 7102 9274 7108 9276
rect 7164 9274 7188 9276
rect 7244 9274 7268 9276
rect 7324 9274 7348 9276
rect 7404 9274 7410 9276
rect 7164 9222 7166 9274
rect 7346 9222 7348 9274
rect 7102 9220 7108 9222
rect 7164 9220 7188 9222
rect 7244 9220 7268 9222
rect 7324 9220 7348 9222
rect 7404 9220 7410 9222
rect 7102 9211 7410 9220
rect 7484 8974 7512 9318
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 7576 8430 7604 8910
rect 7668 8906 7696 9982
rect 7840 9930 7892 9936
rect 7762 9820 8070 9829
rect 7762 9818 7768 9820
rect 7824 9818 7848 9820
rect 7904 9818 7928 9820
rect 7984 9818 8008 9820
rect 8064 9818 8070 9820
rect 7824 9766 7826 9818
rect 8006 9766 8008 9818
rect 7762 9764 7768 9766
rect 7824 9764 7848 9766
rect 7904 9764 7928 9766
rect 7984 9764 8008 9766
rect 8064 9764 8070 9766
rect 7762 9755 8070 9764
rect 8220 9654 8248 10202
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8588 9994 8616 10134
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 9722 8340 9862
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8220 8974 8248 9590
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 8312 8838 8340 9658
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8404 8974 8432 9454
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 7762 8732 8070 8741
rect 7762 8730 7768 8732
rect 7824 8730 7848 8732
rect 7904 8730 7928 8732
rect 7984 8730 8008 8732
rect 8064 8730 8070 8732
rect 7824 8678 7826 8730
rect 8006 8678 8008 8730
rect 7762 8676 7768 8678
rect 7824 8676 7848 8678
rect 7904 8676 7928 8678
rect 7984 8676 8008 8678
rect 8064 8676 8070 8678
rect 7762 8667 8070 8676
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 8312 8294 8340 8774
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 7102 8188 7410 8197
rect 7102 8186 7108 8188
rect 7164 8186 7188 8188
rect 7244 8186 7268 8188
rect 7324 8186 7348 8188
rect 7404 8186 7410 8188
rect 7164 8134 7166 8186
rect 7346 8134 7348 8186
rect 7102 8132 7108 8134
rect 7164 8132 7188 8134
rect 7244 8132 7268 8134
rect 7324 8132 7348 8134
rect 7404 8132 7410 8134
rect 7102 8123 7410 8132
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6656 7410 6684 7686
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5170 7032 5226 7041
rect 4344 6996 4396 7002
rect 4448 6990 4568 7018
rect 4344 6938 4396 6944
rect 4540 6934 4568 6990
rect 5170 6967 5226 6976
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 5276 6866 5304 7142
rect 5998 6896 6054 6905
rect 5264 6860 5316 6866
rect 5998 6831 6054 6840
rect 5264 6802 5316 6808
rect 6012 6798 6040 6831
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 5301 6556 5609 6565
rect 5301 6554 5307 6556
rect 5363 6554 5387 6556
rect 5443 6554 5467 6556
rect 5523 6554 5547 6556
rect 5603 6554 5609 6556
rect 5363 6502 5365 6554
rect 5545 6502 5547 6554
rect 5301 6500 5307 6502
rect 5363 6500 5387 6502
rect 5443 6500 5467 6502
rect 5523 6500 5547 6502
rect 5603 6500 5609 6502
rect 5301 6491 5609 6500
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 3344 5574 3372 5714
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 2840 5468 3148 5477
rect 2840 5466 2846 5468
rect 2902 5466 2926 5468
rect 2982 5466 3006 5468
rect 3062 5466 3086 5468
rect 3142 5466 3148 5468
rect 2902 5414 2904 5466
rect 3084 5414 3086 5466
rect 2840 5412 2846 5414
rect 2902 5412 2926 5414
rect 2982 5412 3006 5414
rect 3062 5412 3086 5414
rect 3142 5412 3148 5414
rect 2840 5403 3148 5412
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 846 4992 902 5001
rect 846 4927 902 4936
rect 1780 4078 1808 5102
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2180 4924 2488 4933
rect 2180 4922 2186 4924
rect 2242 4922 2266 4924
rect 2322 4922 2346 4924
rect 2402 4922 2426 4924
rect 2482 4922 2488 4924
rect 2242 4870 2244 4922
rect 2424 4870 2426 4922
rect 2180 4868 2186 4870
rect 2242 4868 2266 4870
rect 2322 4868 2346 4870
rect 2402 4868 2426 4870
rect 2482 4868 2488 4870
rect 2180 4859 2488 4868
rect 2792 4690 2820 4966
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2884 4622 2912 4966
rect 3344 4690 3372 5510
rect 4172 5234 4200 5782
rect 4264 5642 4292 6190
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4448 5778 4476 6054
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 5234 4476 5510
rect 4540 5370 4568 6258
rect 4641 6012 4949 6021
rect 4641 6010 4647 6012
rect 4703 6010 4727 6012
rect 4783 6010 4807 6012
rect 4863 6010 4887 6012
rect 4943 6010 4949 6012
rect 4703 5958 4705 6010
rect 4885 5958 4887 6010
rect 4641 5956 4647 5958
rect 4703 5956 4727 5958
rect 4783 5956 4807 5958
rect 4863 5956 4887 5958
rect 4943 5956 4949 5958
rect 4641 5947 4949 5956
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5301 5468 5609 5477
rect 5301 5466 5307 5468
rect 5363 5466 5387 5468
rect 5443 5466 5467 5468
rect 5523 5466 5547 5468
rect 5603 5466 5609 5468
rect 5363 5414 5365 5466
rect 5545 5414 5547 5466
rect 5301 5412 5307 5414
rect 5363 5412 5387 5414
rect 5443 5412 5467 5414
rect 5523 5412 5547 5414
rect 5603 5412 5609 5414
rect 5301 5403 5609 5412
rect 5644 5370 5672 5578
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4641 4924 4949 4933
rect 4641 4922 4647 4924
rect 4703 4922 4727 4924
rect 4783 4922 4807 4924
rect 4863 4922 4887 4924
rect 4943 4922 4949 4924
rect 4703 4870 4705 4922
rect 4885 4870 4887 4922
rect 4641 4868 4647 4870
rect 4703 4868 4727 4870
rect 4783 4868 4807 4870
rect 4863 4868 4887 4870
rect 4943 4868 4949 4870
rect 4641 4859 4949 4868
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 2148 4214 2176 4422
rect 2840 4380 3148 4389
rect 2840 4378 2846 4380
rect 2902 4378 2926 4380
rect 2982 4378 3006 4380
rect 3062 4378 3086 4380
rect 3142 4378 3148 4380
rect 2902 4326 2904 4378
rect 3084 4326 3086 4378
rect 2840 4324 2846 4326
rect 2902 4324 2926 4326
rect 2982 4324 3006 4326
rect 3062 4324 3086 4326
rect 3142 4324 3148 4326
rect 2840 4315 3148 4324
rect 2136 4208 2188 4214
rect 2136 4150 2188 4156
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1780 3602 1808 4014
rect 2180 3836 2488 3845
rect 2180 3834 2186 3836
rect 2242 3834 2266 3836
rect 2322 3834 2346 3836
rect 2402 3834 2426 3836
rect 2482 3834 2488 3836
rect 2242 3782 2244 3834
rect 2424 3782 2426 3834
rect 2180 3780 2186 3782
rect 2242 3780 2266 3782
rect 2322 3780 2346 3782
rect 2402 3780 2426 3782
rect 2482 3780 2488 3782
rect 2180 3771 2488 3780
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1964 3194 1992 3470
rect 2840 3292 3148 3301
rect 2840 3290 2846 3292
rect 2902 3290 2926 3292
rect 2982 3290 3006 3292
rect 3062 3290 3086 3292
rect 3142 3290 3148 3292
rect 2902 3238 2904 3290
rect 3084 3238 3086 3290
rect 2840 3236 2846 3238
rect 2902 3236 2926 3238
rect 2982 3236 3006 3238
rect 3062 3236 3086 3238
rect 3142 3236 3148 3238
rect 2840 3227 3148 3236
rect 3252 3194 3280 4422
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3344 2990 3372 4626
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 3194 3648 4082
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3712 3466 3740 3878
rect 3804 3738 3832 4014
rect 4356 4010 4384 4558
rect 4632 4282 4660 4558
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4344 4004 4396 4010
rect 4344 3946 4396 3952
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3988 3194 4016 3878
rect 4641 3836 4949 3845
rect 4641 3834 4647 3836
rect 4703 3834 4727 3836
rect 4783 3834 4807 3836
rect 4863 3834 4887 3836
rect 4943 3834 4949 3836
rect 4703 3782 4705 3834
rect 4885 3782 4887 3834
rect 4641 3780 4647 3782
rect 4703 3780 4727 3782
rect 4783 3780 4807 3782
rect 4863 3780 4887 3782
rect 4943 3780 4949 3782
rect 4641 3771 4949 3780
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 2180 2748 2488 2757
rect 2180 2746 2186 2748
rect 2242 2746 2266 2748
rect 2322 2746 2346 2748
rect 2402 2746 2426 2748
rect 2482 2746 2488 2748
rect 2242 2694 2244 2746
rect 2424 2694 2426 2746
rect 2180 2692 2186 2694
rect 2242 2692 2266 2694
rect 2322 2692 2346 2694
rect 2402 2692 2426 2694
rect 2482 2692 2488 2694
rect 2180 2683 2488 2692
rect 3160 2650 3188 2926
rect 4172 2650 4200 3062
rect 4816 3058 4844 3470
rect 5092 3126 5120 4422
rect 5184 4282 5212 4422
rect 5301 4380 5609 4389
rect 5301 4378 5307 4380
rect 5363 4378 5387 4380
rect 5443 4378 5467 4380
rect 5523 4378 5547 4380
rect 5603 4378 5609 4380
rect 5363 4326 5365 4378
rect 5545 4326 5547 4378
rect 5301 4324 5307 4326
rect 5363 4324 5387 4326
rect 5443 4324 5467 4326
rect 5523 4324 5547 4326
rect 5603 4324 5609 4326
rect 5301 4315 5609 4324
rect 5644 4282 5672 4558
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4641 2748 4949 2757
rect 4641 2746 4647 2748
rect 4703 2746 4727 2748
rect 4783 2746 4807 2748
rect 4863 2746 4887 2748
rect 4943 2746 4949 2748
rect 4703 2694 4705 2746
rect 4885 2694 4887 2746
rect 4641 2692 4647 2694
rect 4703 2692 4727 2694
rect 4783 2692 4807 2694
rect 4863 2692 4887 2694
rect 4943 2692 4949 2694
rect 4641 2683 4949 2692
rect 5184 2650 5212 4014
rect 5301 3292 5609 3301
rect 5301 3290 5307 3292
rect 5363 3290 5387 3292
rect 5443 3290 5467 3292
rect 5523 3290 5547 3292
rect 5603 3290 5609 3292
rect 5363 3238 5365 3290
rect 5545 3238 5547 3290
rect 5301 3236 5307 3238
rect 5363 3236 5387 3238
rect 5443 3236 5467 3238
rect 5523 3236 5547 3238
rect 5603 3236 5609 3238
rect 5301 3227 5609 3236
rect 5644 3194 5672 4014
rect 5736 3466 5764 4694
rect 6104 4690 6132 5646
rect 6196 5574 6224 6666
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6458 6316 6598
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6380 6322 6408 7278
rect 7102 7100 7410 7109
rect 7102 7098 7108 7100
rect 7164 7098 7188 7100
rect 7244 7098 7268 7100
rect 7324 7098 7348 7100
rect 7404 7098 7410 7100
rect 7164 7046 7166 7098
rect 7346 7046 7348 7098
rect 7102 7044 7108 7046
rect 7164 7044 7188 7046
rect 7244 7044 7268 7046
rect 7324 7044 7348 7046
rect 7404 7044 7410 7046
rect 7102 7035 7410 7044
rect 7576 7002 7604 7822
rect 7762 7644 8070 7653
rect 7762 7642 7768 7644
rect 7824 7642 7848 7644
rect 7904 7642 7928 7644
rect 7984 7642 8008 7644
rect 8064 7642 8070 7644
rect 7824 7590 7826 7642
rect 8006 7590 8008 7642
rect 7762 7588 7768 7590
rect 7824 7588 7848 7590
rect 7904 7588 7928 7590
rect 7984 7588 8008 7590
rect 8064 7588 8070 7590
rect 7762 7579 8070 7588
rect 8128 7478 8156 7822
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7286 6896 7342 6905
rect 8312 6866 8340 7686
rect 8588 7274 8616 9930
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 9042 9076 9318
rect 9232 9178 9260 9930
rect 10223 9820 10531 9829
rect 10223 9818 10229 9820
rect 10285 9818 10309 9820
rect 10365 9818 10389 9820
rect 10445 9818 10469 9820
rect 10525 9818 10531 9820
rect 10285 9766 10287 9818
rect 10467 9766 10469 9818
rect 10223 9764 10229 9766
rect 10285 9764 10309 9766
rect 10365 9764 10389 9766
rect 10445 9764 10469 9766
rect 10525 9764 10531 9766
rect 10223 9755 10531 9764
rect 10612 9625 10640 9998
rect 10598 9616 10654 9625
rect 10704 9586 10732 10066
rect 10598 9551 10654 9560
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 9563 9276 9871 9285
rect 9563 9274 9569 9276
rect 9625 9274 9649 9276
rect 9705 9274 9729 9276
rect 9785 9274 9809 9276
rect 9865 9274 9871 9276
rect 9625 9222 9627 9274
rect 9807 9222 9809 9274
rect 9563 9220 9569 9222
rect 9625 9220 9649 9222
rect 9705 9220 9729 9222
rect 9785 9220 9809 9222
rect 9865 9220 9871 9222
rect 9563 9211 9871 9220
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 10598 8936 10654 8945
rect 10598 8871 10654 8880
rect 10223 8732 10531 8741
rect 10223 8730 10229 8732
rect 10285 8730 10309 8732
rect 10365 8730 10389 8732
rect 10445 8730 10469 8732
rect 10525 8730 10531 8732
rect 10285 8678 10287 8730
rect 10467 8678 10469 8730
rect 10223 8676 10229 8678
rect 10285 8676 10309 8678
rect 10365 8676 10389 8678
rect 10445 8676 10469 8678
rect 10525 8676 10531 8678
rect 10223 8667 10531 8676
rect 10612 8634 10640 8871
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 7286 6831 7342 6840
rect 8300 6860 8352 6866
rect 7300 6662 7328 6831
rect 8300 6802 8352 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6460 6316 6512 6322
rect 6564 6304 6592 6394
rect 6656 6322 6684 6598
rect 7300 6390 7328 6598
rect 7762 6556 8070 6565
rect 7762 6554 7768 6556
rect 7824 6554 7848 6556
rect 7904 6554 7928 6556
rect 7984 6554 8008 6556
rect 8064 6554 8070 6556
rect 7824 6502 7826 6554
rect 8006 6502 8008 6554
rect 7762 6500 7768 6502
rect 7824 6500 7848 6502
rect 7904 6500 7928 6502
rect 7984 6500 8008 6502
rect 8064 6500 8070 6502
rect 7762 6491 8070 6500
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 6512 6276 6592 6304
rect 6644 6316 6696 6322
rect 6460 6258 6512 6264
rect 6644 6258 6696 6264
rect 6380 5914 6408 6258
rect 7024 5914 7052 6326
rect 7102 6012 7410 6021
rect 7102 6010 7108 6012
rect 7164 6010 7188 6012
rect 7244 6010 7268 6012
rect 7324 6010 7348 6012
rect 7404 6010 7410 6012
rect 7164 5958 7166 6010
rect 7346 5958 7348 6010
rect 7102 5956 7108 5958
rect 7164 5956 7188 5958
rect 7244 5956 7268 5958
rect 7324 5956 7348 5958
rect 7404 5956 7410 5958
rect 7102 5947 7410 5956
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 8312 5778 8340 6598
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8404 5642 8432 6394
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6196 5234 6224 5510
rect 6380 5370 6408 5578
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 4826 6776 5170
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6932 4690 6960 4966
rect 7102 4924 7410 4933
rect 7102 4922 7108 4924
rect 7164 4922 7188 4924
rect 7244 4922 7268 4924
rect 7324 4922 7348 4924
rect 7404 4922 7410 4924
rect 7164 4870 7166 4922
rect 7346 4870 7348 4922
rect 7102 4868 7108 4870
rect 7164 4868 7188 4870
rect 7244 4868 7268 4870
rect 7324 4868 7348 4870
rect 7404 4868 7410 4870
rect 7102 4859 7410 4868
rect 7576 4826 7604 5510
rect 7668 4826 7696 5510
rect 7762 5468 8070 5477
rect 7762 5466 7768 5468
rect 7824 5466 7848 5468
rect 7904 5466 7928 5468
rect 7984 5466 8008 5468
rect 8064 5466 8070 5468
rect 7824 5414 7826 5466
rect 8006 5414 8008 5466
rect 7762 5412 7768 5414
rect 7824 5412 7848 5414
rect 7904 5412 7928 5414
rect 7984 5412 8008 5414
rect 8064 5412 8070 5414
rect 7762 5403 8070 5412
rect 8312 5234 8340 5578
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8220 4826 8248 5170
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5828 3738 5856 4558
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 6104 2650 6132 4014
rect 6288 2650 6316 4422
rect 7762 4380 8070 4389
rect 7762 4378 7768 4380
rect 7824 4378 7848 4380
rect 7904 4378 7928 4380
rect 7984 4378 8008 4380
rect 8064 4378 8070 4380
rect 7824 4326 7826 4378
rect 8006 4326 8008 4378
rect 7762 4324 7768 4326
rect 7824 4324 7848 4326
rect 7904 4324 7928 4326
rect 7984 4324 8008 4326
rect 8064 4324 8070 4326
rect 7762 4315 8070 4324
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 6920 4004 6972 4010
rect 6920 3946 6972 3952
rect 6932 3058 6960 3946
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 7024 3194 7052 3878
rect 7102 3836 7410 3845
rect 7102 3834 7108 3836
rect 7164 3834 7188 3836
rect 7244 3834 7268 3836
rect 7324 3834 7348 3836
rect 7404 3834 7410 3836
rect 7164 3782 7166 3834
rect 7346 3782 7348 3834
rect 7102 3780 7108 3782
rect 7164 3780 7188 3782
rect 7244 3780 7268 3782
rect 7324 3780 7348 3782
rect 7404 3780 7410 3782
rect 7102 3771 7410 3780
rect 7576 3738 7604 4014
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 8312 3534 8340 5170
rect 8496 4690 8524 6054
rect 8588 5846 8616 6734
rect 8680 6662 8708 7278
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8772 5914 8800 7482
rect 9140 7410 9168 8230
rect 9563 8188 9871 8197
rect 9563 8186 9569 8188
rect 9625 8186 9649 8188
rect 9705 8186 9729 8188
rect 9785 8186 9809 8188
rect 9865 8186 9871 8188
rect 9625 8134 9627 8186
rect 9807 8134 9809 8186
rect 9563 8132 9569 8134
rect 9625 8132 9649 8134
rect 9705 8132 9729 8134
rect 9785 8132 9809 8134
rect 9865 8132 9871 8134
rect 9563 8123 9871 8132
rect 9968 7546 9996 8434
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 9956 7540 10008 7546
rect 9956 7482 10008 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8864 5914 8892 7278
rect 8956 6118 8984 7278
rect 9563 7100 9871 7109
rect 9563 7098 9569 7100
rect 9625 7098 9649 7100
rect 9705 7098 9729 7100
rect 9785 7098 9809 7100
rect 9865 7098 9871 7100
rect 9625 7046 9627 7098
rect 9807 7046 9809 7098
rect 9563 7044 9569 7046
rect 9625 7044 9649 7046
rect 9705 7044 9729 7046
rect 9785 7044 9809 7046
rect 9865 7044 9871 7046
rect 9563 7035 9871 7044
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9600 6254 9628 6734
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8588 5166 8616 5782
rect 8864 5370 8892 5850
rect 9324 5710 9352 6190
rect 9563 6012 9871 6021
rect 9563 6010 9569 6012
rect 9625 6010 9649 6012
rect 9705 6010 9729 6012
rect 9785 6010 9809 6012
rect 9865 6010 9871 6012
rect 9625 5958 9627 6010
rect 9807 5958 9809 6010
rect 9563 5956 9569 5958
rect 9625 5956 9649 5958
rect 9705 5956 9729 5958
rect 9785 5956 9809 5958
rect 9865 5956 9871 5958
rect 9563 5947 9871 5956
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 9324 5234 9352 5646
rect 10152 5370 10180 7822
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10223 7644 10531 7653
rect 10223 7642 10229 7644
rect 10285 7642 10309 7644
rect 10365 7642 10389 7644
rect 10445 7642 10469 7644
rect 10525 7642 10531 7644
rect 10285 7590 10287 7642
rect 10467 7590 10469 7642
rect 10223 7588 10229 7590
rect 10285 7588 10309 7590
rect 10365 7588 10389 7590
rect 10445 7588 10469 7590
rect 10525 7588 10531 7590
rect 10223 7579 10531 7588
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 6798 10640 7142
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10223 6556 10531 6565
rect 10223 6554 10229 6556
rect 10285 6554 10309 6556
rect 10365 6554 10389 6556
rect 10445 6554 10469 6556
rect 10525 6554 10531 6556
rect 10285 6502 10287 6554
rect 10467 6502 10469 6554
rect 10223 6500 10229 6502
rect 10285 6500 10309 6502
rect 10365 6500 10389 6502
rect 10445 6500 10469 6502
rect 10525 6500 10531 6502
rect 10223 6491 10531 6500
rect 10704 6322 10732 7686
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5642 10456 6054
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10223 5468 10531 5477
rect 10223 5466 10229 5468
rect 10285 5466 10309 5468
rect 10365 5466 10389 5468
rect 10445 5466 10469 5468
rect 10525 5466 10531 5468
rect 10285 5414 10287 5466
rect 10467 5414 10469 5466
rect 10223 5412 10229 5414
rect 10285 5412 10309 5414
rect 10365 5412 10389 5414
rect 10445 5412 10469 5414
rect 10525 5412 10531 5414
rect 10223 5403 10531 5412
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8680 4622 8708 5034
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8864 4078 8892 4966
rect 9324 4826 9352 5170
rect 9563 4924 9871 4933
rect 9563 4922 9569 4924
rect 9625 4922 9649 4924
rect 9705 4922 9729 4924
rect 9785 4922 9809 4924
rect 9865 4922 9871 4924
rect 9625 4870 9627 4922
rect 9807 4870 9809 4922
rect 9563 4868 9569 4870
rect 9625 4868 9649 4870
rect 9705 4868 9729 4870
rect 9785 4868 9809 4870
rect 9865 4868 9871 4870
rect 9563 4859 9871 4868
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9600 4282 9628 4490
rect 10060 4282 10088 5170
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10336 4826 10364 5102
rect 10598 4856 10654 4865
rect 10324 4820 10376 4826
rect 10598 4791 10654 4800
rect 10324 4762 10376 4768
rect 10612 4622 10640 4791
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 3194 7696 3402
rect 7762 3292 8070 3301
rect 7762 3290 7768 3292
rect 7824 3290 7848 3292
rect 7904 3290 7928 3292
rect 7984 3290 8008 3292
rect 8064 3290 8070 3292
rect 7824 3238 7826 3290
rect 8006 3238 8008 3290
rect 7762 3236 7768 3238
rect 7824 3236 7848 3238
rect 7904 3236 7928 3238
rect 7984 3236 8008 3238
rect 8064 3236 8070 3238
rect 7762 3227 8070 3236
rect 8312 3194 8340 3470
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8404 3126 8432 3334
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7104 2984 7156 2990
rect 7024 2932 7104 2938
rect 7024 2926 7156 2932
rect 7024 2910 7144 2926
rect 7024 2650 7052 2910
rect 7102 2748 7410 2757
rect 7102 2746 7108 2748
rect 7164 2746 7188 2748
rect 7244 2746 7268 2748
rect 7324 2746 7348 2748
rect 7404 2746 7410 2748
rect 7164 2694 7166 2746
rect 7346 2694 7348 2746
rect 7102 2692 7108 2694
rect 7164 2692 7188 2694
rect 7244 2692 7268 2694
rect 7324 2692 7348 2694
rect 7404 2692 7410 2694
rect 7102 2683 7410 2692
rect 8496 2650 8524 4014
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 3534 8616 3878
rect 8956 3738 8984 4082
rect 9563 3836 9871 3845
rect 9563 3834 9569 3836
rect 9625 3834 9649 3836
rect 9705 3834 9729 3836
rect 9785 3834 9809 3836
rect 9865 3834 9871 3836
rect 9625 3782 9627 3834
rect 9807 3782 9809 3834
rect 9563 3780 9569 3782
rect 9625 3780 9649 3782
rect 9705 3780 9729 3782
rect 9785 3780 9809 3782
rect 9865 3780 9871 3782
rect 9563 3771 9871 3780
rect 9968 3738 9996 4150
rect 10152 4146 10180 4422
rect 10223 4380 10531 4389
rect 10223 4378 10229 4380
rect 10285 4378 10309 4380
rect 10365 4378 10389 4380
rect 10445 4378 10469 4380
rect 10525 4378 10531 4380
rect 10285 4326 10287 4378
rect 10467 4326 10469 4378
rect 10223 4324 10229 4326
rect 10285 4324 10309 4326
rect 10365 4324 10389 4326
rect 10445 4324 10469 4326
rect 10525 4324 10531 4326
rect 10223 4315 10531 4324
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3738 10456 3878
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 9588 3528 9640 3534
rect 10600 3528 10652 3534
rect 9588 3470 9640 3476
rect 10598 3496 10600 3505
rect 10652 3496 10654 3505
rect 9600 3194 9628 3470
rect 10598 3431 10654 3440
rect 10223 3292 10531 3301
rect 10223 3290 10229 3292
rect 10285 3290 10309 3292
rect 10365 3290 10389 3292
rect 10445 3290 10469 3292
rect 10525 3290 10531 3292
rect 10285 3238 10287 3290
rect 10467 3238 10469 3290
rect 10223 3236 10229 3238
rect 10285 3236 10309 3238
rect 10365 3236 10389 3238
rect 10445 3236 10469 3238
rect 10525 3236 10531 3238
rect 10223 3227 10531 3236
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9563 2748 9871 2757
rect 9563 2746 9569 2748
rect 9625 2746 9649 2748
rect 9705 2746 9729 2748
rect 9785 2746 9809 2748
rect 9865 2746 9871 2748
rect 9625 2694 9627 2746
rect 9807 2694 9809 2746
rect 9563 2692 9569 2694
rect 9625 2692 9649 2694
rect 9705 2692 9729 2694
rect 9785 2692 9809 2694
rect 9865 2692 9871 2694
rect 9563 2683 9871 2692
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 2840 2204 3148 2213
rect 2840 2202 2846 2204
rect 2902 2202 2926 2204
rect 2982 2202 3006 2204
rect 3062 2202 3086 2204
rect 3142 2202 3148 2204
rect 2902 2150 2904 2202
rect 3084 2150 3086 2202
rect 2840 2148 2846 2150
rect 2902 2148 2926 2150
rect 2982 2148 3006 2150
rect 3062 2148 3086 2150
rect 3142 2148 3148 2150
rect 2840 2139 3148 2148
rect 3252 800 3280 2382
rect 3896 800 3924 2382
rect 5184 800 5212 2382
rect 5301 2204 5609 2213
rect 5301 2202 5307 2204
rect 5363 2202 5387 2204
rect 5443 2202 5467 2204
rect 5523 2202 5547 2204
rect 5603 2202 5609 2204
rect 5363 2150 5365 2202
rect 5545 2150 5547 2202
rect 5301 2148 5307 2150
rect 5363 2148 5387 2150
rect 5443 2148 5467 2150
rect 5523 2148 5547 2150
rect 5603 2148 5609 2150
rect 5301 2139 5609 2148
rect 5828 800 5856 2382
rect 6472 800 6500 2382
rect 7116 800 7144 2382
rect 7762 2204 8070 2213
rect 7762 2202 7768 2204
rect 7824 2202 7848 2204
rect 7904 2202 7928 2204
rect 7984 2202 8008 2204
rect 8064 2202 8070 2204
rect 7824 2150 7826 2202
rect 8006 2150 8008 2202
rect 7762 2148 7768 2150
rect 7824 2148 7848 2150
rect 7904 2148 7928 2150
rect 7984 2148 8008 2150
rect 8064 2148 8070 2150
rect 7762 2139 8070 2148
rect 8404 800 8432 2382
rect 10223 2204 10531 2213
rect 10223 2202 10229 2204
rect 10285 2202 10309 2204
rect 10365 2202 10389 2204
rect 10445 2202 10469 2204
rect 10525 2202 10531 2204
rect 10285 2150 10287 2202
rect 10467 2150 10469 2202
rect 10223 2148 10229 2150
rect 10285 2148 10309 2150
rect 10365 2148 10389 2150
rect 10445 2148 10469 2150
rect 10525 2148 10531 2150
rect 10223 2139 10531 2148
rect 18 0 74 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 8390 0 8446 800
<< via2 >>
rect 2846 11994 2902 11996
rect 2926 11994 2982 11996
rect 3006 11994 3062 11996
rect 3086 11994 3142 11996
rect 2846 11942 2892 11994
rect 2892 11942 2902 11994
rect 2926 11942 2956 11994
rect 2956 11942 2968 11994
rect 2968 11942 2982 11994
rect 3006 11942 3020 11994
rect 3020 11942 3032 11994
rect 3032 11942 3062 11994
rect 3086 11942 3096 11994
rect 3096 11942 3142 11994
rect 2846 11940 2902 11942
rect 2926 11940 2982 11942
rect 3006 11940 3062 11942
rect 3086 11940 3142 11942
rect 5307 11994 5363 11996
rect 5387 11994 5443 11996
rect 5467 11994 5523 11996
rect 5547 11994 5603 11996
rect 5307 11942 5353 11994
rect 5353 11942 5363 11994
rect 5387 11942 5417 11994
rect 5417 11942 5429 11994
rect 5429 11942 5443 11994
rect 5467 11942 5481 11994
rect 5481 11942 5493 11994
rect 5493 11942 5523 11994
rect 5547 11942 5557 11994
rect 5557 11942 5603 11994
rect 5307 11940 5363 11942
rect 5387 11940 5443 11942
rect 5467 11940 5523 11942
rect 5547 11940 5603 11942
rect 7768 11994 7824 11996
rect 7848 11994 7904 11996
rect 7928 11994 7984 11996
rect 8008 11994 8064 11996
rect 7768 11942 7814 11994
rect 7814 11942 7824 11994
rect 7848 11942 7878 11994
rect 7878 11942 7890 11994
rect 7890 11942 7904 11994
rect 7928 11942 7942 11994
rect 7942 11942 7954 11994
rect 7954 11942 7984 11994
rect 8008 11942 8018 11994
rect 8018 11942 8064 11994
rect 7768 11940 7824 11942
rect 7848 11940 7904 11942
rect 7928 11940 7984 11942
rect 8008 11940 8064 11942
rect 10229 11994 10285 11996
rect 10309 11994 10365 11996
rect 10389 11994 10445 11996
rect 10469 11994 10525 11996
rect 10229 11942 10275 11994
rect 10275 11942 10285 11994
rect 10309 11942 10339 11994
rect 10339 11942 10351 11994
rect 10351 11942 10365 11994
rect 10389 11942 10403 11994
rect 10403 11942 10415 11994
rect 10415 11942 10445 11994
rect 10469 11942 10479 11994
rect 10479 11942 10525 11994
rect 10229 11940 10285 11942
rect 10309 11940 10365 11942
rect 10389 11940 10445 11942
rect 10469 11940 10525 11942
rect 2186 11450 2242 11452
rect 2266 11450 2322 11452
rect 2346 11450 2402 11452
rect 2426 11450 2482 11452
rect 2186 11398 2232 11450
rect 2232 11398 2242 11450
rect 2266 11398 2296 11450
rect 2296 11398 2308 11450
rect 2308 11398 2322 11450
rect 2346 11398 2360 11450
rect 2360 11398 2372 11450
rect 2372 11398 2402 11450
rect 2426 11398 2436 11450
rect 2436 11398 2482 11450
rect 2186 11396 2242 11398
rect 2266 11396 2322 11398
rect 2346 11396 2402 11398
rect 2426 11396 2482 11398
rect 846 10376 902 10432
rect 2186 10362 2242 10364
rect 2266 10362 2322 10364
rect 2346 10362 2402 10364
rect 2426 10362 2482 10364
rect 2186 10310 2232 10362
rect 2232 10310 2242 10362
rect 2266 10310 2296 10362
rect 2296 10310 2308 10362
rect 2308 10310 2322 10362
rect 2346 10310 2360 10362
rect 2360 10310 2372 10362
rect 2372 10310 2402 10362
rect 2426 10310 2436 10362
rect 2436 10310 2482 10362
rect 2186 10308 2242 10310
rect 2266 10308 2322 10310
rect 2346 10308 2402 10310
rect 2426 10308 2482 10310
rect 2846 10906 2902 10908
rect 2926 10906 2982 10908
rect 3006 10906 3062 10908
rect 3086 10906 3142 10908
rect 2846 10854 2892 10906
rect 2892 10854 2902 10906
rect 2926 10854 2956 10906
rect 2956 10854 2968 10906
rect 2968 10854 2982 10906
rect 3006 10854 3020 10906
rect 3020 10854 3032 10906
rect 3032 10854 3062 10906
rect 3086 10854 3096 10906
rect 3096 10854 3142 10906
rect 2846 10852 2902 10854
rect 2926 10852 2982 10854
rect 3006 10852 3062 10854
rect 3086 10852 3142 10854
rect 1398 8200 1454 8256
rect 2186 9274 2242 9276
rect 2266 9274 2322 9276
rect 2346 9274 2402 9276
rect 2426 9274 2482 9276
rect 2186 9222 2232 9274
rect 2232 9222 2242 9274
rect 2266 9222 2296 9274
rect 2296 9222 2308 9274
rect 2308 9222 2322 9274
rect 2346 9222 2360 9274
rect 2360 9222 2372 9274
rect 2372 9222 2402 9274
rect 2426 9222 2436 9274
rect 2436 9222 2482 9274
rect 2186 9220 2242 9222
rect 2266 9220 2322 9222
rect 2346 9220 2402 9222
rect 2426 9220 2482 9222
rect 2846 9818 2902 9820
rect 2926 9818 2982 9820
rect 3006 9818 3062 9820
rect 3086 9818 3142 9820
rect 2846 9766 2892 9818
rect 2892 9766 2902 9818
rect 2926 9766 2956 9818
rect 2956 9766 2968 9818
rect 2968 9766 2982 9818
rect 3006 9766 3020 9818
rect 3020 9766 3032 9818
rect 3032 9766 3062 9818
rect 3086 9766 3096 9818
rect 3096 9766 3142 9818
rect 2846 9764 2902 9766
rect 2926 9764 2982 9766
rect 3006 9764 3062 9766
rect 3086 9764 3142 9766
rect 2846 8730 2902 8732
rect 2926 8730 2982 8732
rect 3006 8730 3062 8732
rect 3086 8730 3142 8732
rect 2846 8678 2892 8730
rect 2892 8678 2902 8730
rect 2926 8678 2956 8730
rect 2956 8678 2968 8730
rect 2968 8678 2982 8730
rect 3006 8678 3020 8730
rect 3020 8678 3032 8730
rect 3032 8678 3062 8730
rect 3086 8678 3096 8730
rect 3096 8678 3142 8730
rect 2846 8676 2902 8678
rect 2926 8676 2982 8678
rect 3006 8676 3062 8678
rect 3086 8676 3142 8678
rect 2186 8186 2242 8188
rect 2266 8186 2322 8188
rect 2346 8186 2402 8188
rect 2426 8186 2482 8188
rect 2186 8134 2232 8186
rect 2232 8134 2242 8186
rect 2266 8134 2296 8186
rect 2296 8134 2308 8186
rect 2308 8134 2322 8186
rect 2346 8134 2360 8186
rect 2360 8134 2372 8186
rect 2372 8134 2402 8186
rect 2426 8134 2436 8186
rect 2436 8134 2482 8186
rect 2186 8132 2242 8134
rect 2266 8132 2322 8134
rect 2346 8132 2402 8134
rect 2426 8132 2482 8134
rect 846 7656 902 7712
rect 2846 7642 2902 7644
rect 2926 7642 2982 7644
rect 3006 7642 3062 7644
rect 3086 7642 3142 7644
rect 2846 7590 2892 7642
rect 2892 7590 2902 7642
rect 2926 7590 2956 7642
rect 2956 7590 2968 7642
rect 2968 7590 2982 7642
rect 3006 7590 3020 7642
rect 3020 7590 3032 7642
rect 3032 7590 3062 7642
rect 3086 7590 3096 7642
rect 3096 7590 3142 7642
rect 2846 7588 2902 7590
rect 2926 7588 2982 7590
rect 3006 7588 3062 7590
rect 3086 7588 3142 7590
rect 2186 7098 2242 7100
rect 2266 7098 2322 7100
rect 2346 7098 2402 7100
rect 2426 7098 2482 7100
rect 2186 7046 2232 7098
rect 2232 7046 2242 7098
rect 2266 7046 2296 7098
rect 2296 7046 2308 7098
rect 2308 7046 2322 7098
rect 2346 7046 2360 7098
rect 2360 7046 2372 7098
rect 2372 7046 2402 7098
rect 2426 7046 2436 7098
rect 2436 7046 2482 7098
rect 2186 7044 2242 7046
rect 2266 7044 2322 7046
rect 2346 7044 2402 7046
rect 2426 7044 2482 7046
rect 1398 6840 1454 6896
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 4647 11450 4703 11452
rect 4727 11450 4783 11452
rect 4807 11450 4863 11452
rect 4887 11450 4943 11452
rect 4647 11398 4693 11450
rect 4693 11398 4703 11450
rect 4727 11398 4757 11450
rect 4757 11398 4769 11450
rect 4769 11398 4783 11450
rect 4807 11398 4821 11450
rect 4821 11398 4833 11450
rect 4833 11398 4863 11450
rect 4887 11398 4897 11450
rect 4897 11398 4943 11450
rect 4647 11396 4703 11398
rect 4727 11396 4783 11398
rect 4807 11396 4863 11398
rect 4887 11396 4943 11398
rect 7108 11450 7164 11452
rect 7188 11450 7244 11452
rect 7268 11450 7324 11452
rect 7348 11450 7404 11452
rect 7108 11398 7154 11450
rect 7154 11398 7164 11450
rect 7188 11398 7218 11450
rect 7218 11398 7230 11450
rect 7230 11398 7244 11450
rect 7268 11398 7282 11450
rect 7282 11398 7294 11450
rect 7294 11398 7324 11450
rect 7348 11398 7358 11450
rect 7358 11398 7404 11450
rect 7108 11396 7164 11398
rect 7188 11396 7244 11398
rect 7268 11396 7324 11398
rect 7348 11396 7404 11398
rect 9569 11450 9625 11452
rect 9649 11450 9705 11452
rect 9729 11450 9785 11452
rect 9809 11450 9865 11452
rect 9569 11398 9615 11450
rect 9615 11398 9625 11450
rect 9649 11398 9679 11450
rect 9679 11398 9691 11450
rect 9691 11398 9705 11450
rect 9729 11398 9743 11450
rect 9743 11398 9755 11450
rect 9755 11398 9785 11450
rect 9809 11398 9819 11450
rect 9819 11398 9865 11450
rect 9569 11396 9625 11398
rect 9649 11396 9705 11398
rect 9729 11396 9785 11398
rect 9809 11396 9865 11398
rect 5307 10906 5363 10908
rect 5387 10906 5443 10908
rect 5467 10906 5523 10908
rect 5547 10906 5603 10908
rect 5307 10854 5353 10906
rect 5353 10854 5363 10906
rect 5387 10854 5417 10906
rect 5417 10854 5429 10906
rect 5429 10854 5443 10906
rect 5467 10854 5481 10906
rect 5481 10854 5493 10906
rect 5493 10854 5523 10906
rect 5547 10854 5557 10906
rect 5557 10854 5603 10906
rect 5307 10852 5363 10854
rect 5387 10852 5443 10854
rect 5467 10852 5523 10854
rect 5547 10852 5603 10854
rect 4647 10362 4703 10364
rect 4727 10362 4783 10364
rect 4807 10362 4863 10364
rect 4887 10362 4943 10364
rect 4647 10310 4693 10362
rect 4693 10310 4703 10362
rect 4727 10310 4757 10362
rect 4757 10310 4769 10362
rect 4769 10310 4783 10362
rect 4807 10310 4821 10362
rect 4821 10310 4833 10362
rect 4833 10310 4863 10362
rect 4887 10310 4897 10362
rect 4897 10310 4943 10362
rect 4647 10308 4703 10310
rect 4727 10308 4783 10310
rect 4807 10308 4863 10310
rect 4887 10308 4943 10310
rect 7108 10362 7164 10364
rect 7188 10362 7244 10364
rect 7268 10362 7324 10364
rect 7348 10362 7404 10364
rect 7108 10310 7154 10362
rect 7154 10310 7164 10362
rect 7188 10310 7218 10362
rect 7218 10310 7230 10362
rect 7230 10310 7244 10362
rect 7268 10310 7282 10362
rect 7282 10310 7294 10362
rect 7294 10310 7324 10362
rect 7348 10310 7358 10362
rect 7358 10310 7404 10362
rect 7108 10308 7164 10310
rect 7188 10308 7244 10310
rect 7268 10308 7324 10310
rect 7348 10308 7404 10310
rect 7768 10906 7824 10908
rect 7848 10906 7904 10908
rect 7928 10906 7984 10908
rect 8008 10906 8064 10908
rect 7768 10854 7814 10906
rect 7814 10854 7824 10906
rect 7848 10854 7878 10906
rect 7878 10854 7890 10906
rect 7890 10854 7904 10906
rect 7928 10854 7942 10906
rect 7942 10854 7954 10906
rect 7954 10854 7984 10906
rect 8008 10854 8018 10906
rect 8018 10854 8064 10906
rect 7768 10852 7824 10854
rect 7848 10852 7904 10854
rect 7928 10852 7984 10854
rect 8008 10852 8064 10854
rect 5307 9818 5363 9820
rect 5387 9818 5443 9820
rect 5467 9818 5523 9820
rect 5547 9818 5603 9820
rect 5307 9766 5353 9818
rect 5353 9766 5363 9818
rect 5387 9766 5417 9818
rect 5417 9766 5429 9818
rect 5429 9766 5443 9818
rect 5467 9766 5481 9818
rect 5481 9766 5493 9818
rect 5493 9766 5523 9818
rect 5547 9766 5557 9818
rect 5557 9766 5603 9818
rect 5307 9764 5363 9766
rect 5387 9764 5443 9766
rect 5467 9764 5523 9766
rect 5547 9764 5603 9766
rect 4647 9274 4703 9276
rect 4727 9274 4783 9276
rect 4807 9274 4863 9276
rect 4887 9274 4943 9276
rect 4647 9222 4693 9274
rect 4693 9222 4703 9274
rect 4727 9222 4757 9274
rect 4757 9222 4769 9274
rect 4769 9222 4783 9274
rect 4807 9222 4821 9274
rect 4821 9222 4833 9274
rect 4833 9222 4863 9274
rect 4887 9222 4897 9274
rect 4897 9222 4943 9274
rect 4647 9220 4703 9222
rect 4727 9220 4783 9222
rect 4807 9220 4863 9222
rect 4887 9220 4943 9222
rect 2846 6554 2902 6556
rect 2926 6554 2982 6556
rect 3006 6554 3062 6556
rect 3086 6554 3142 6556
rect 2846 6502 2892 6554
rect 2892 6502 2902 6554
rect 2926 6502 2956 6554
rect 2956 6502 2968 6554
rect 2968 6502 2982 6554
rect 3006 6502 3020 6554
rect 3020 6502 3032 6554
rect 3032 6502 3062 6554
rect 3086 6502 3096 6554
rect 3096 6502 3142 6554
rect 2846 6500 2902 6502
rect 2926 6500 2982 6502
rect 3006 6500 3062 6502
rect 3086 6500 3142 6502
rect 1398 5480 1454 5536
rect 2186 6010 2242 6012
rect 2266 6010 2322 6012
rect 2346 6010 2402 6012
rect 2426 6010 2482 6012
rect 2186 5958 2232 6010
rect 2232 5958 2242 6010
rect 2266 5958 2296 6010
rect 2296 5958 2308 6010
rect 2308 5958 2322 6010
rect 2346 5958 2360 6010
rect 2360 5958 2372 6010
rect 2372 5958 2402 6010
rect 2426 5958 2436 6010
rect 2436 5958 2482 6010
rect 2186 5956 2242 5958
rect 2266 5956 2322 5958
rect 2346 5956 2402 5958
rect 2426 5956 2482 5958
rect 5307 8730 5363 8732
rect 5387 8730 5443 8732
rect 5467 8730 5523 8732
rect 5547 8730 5603 8732
rect 5307 8678 5353 8730
rect 5353 8678 5363 8730
rect 5387 8678 5417 8730
rect 5417 8678 5429 8730
rect 5429 8678 5443 8730
rect 5467 8678 5481 8730
rect 5481 8678 5493 8730
rect 5493 8678 5523 8730
rect 5547 8678 5557 8730
rect 5557 8678 5603 8730
rect 5307 8676 5363 8678
rect 5387 8676 5443 8678
rect 5467 8676 5523 8678
rect 5547 8676 5603 8678
rect 4647 8186 4703 8188
rect 4727 8186 4783 8188
rect 4807 8186 4863 8188
rect 4887 8186 4943 8188
rect 4647 8134 4693 8186
rect 4693 8134 4703 8186
rect 4727 8134 4757 8186
rect 4757 8134 4769 8186
rect 4769 8134 4783 8186
rect 4807 8134 4821 8186
rect 4821 8134 4833 8186
rect 4833 8134 4863 8186
rect 4887 8134 4897 8186
rect 4897 8134 4943 8186
rect 4647 8132 4703 8134
rect 4727 8132 4783 8134
rect 4807 8132 4863 8134
rect 4887 8132 4943 8134
rect 5307 7642 5363 7644
rect 5387 7642 5443 7644
rect 5467 7642 5523 7644
rect 5547 7642 5603 7644
rect 5307 7590 5353 7642
rect 5353 7590 5363 7642
rect 5387 7590 5417 7642
rect 5417 7590 5429 7642
rect 5429 7590 5443 7642
rect 5467 7590 5481 7642
rect 5481 7590 5493 7642
rect 5493 7590 5523 7642
rect 5547 7590 5557 7642
rect 5557 7590 5603 7642
rect 5307 7588 5363 7590
rect 5387 7588 5443 7590
rect 5467 7588 5523 7590
rect 5547 7588 5603 7590
rect 4647 7098 4703 7100
rect 4727 7098 4783 7100
rect 4807 7098 4863 7100
rect 4887 7098 4943 7100
rect 4647 7046 4693 7098
rect 4693 7046 4703 7098
rect 4727 7046 4757 7098
rect 4757 7046 4769 7098
rect 4769 7046 4783 7098
rect 4807 7046 4821 7098
rect 4821 7046 4833 7098
rect 4833 7046 4863 7098
rect 4887 7046 4897 7098
rect 4897 7046 4943 7098
rect 4647 7044 4703 7046
rect 4727 7044 4783 7046
rect 4807 7044 4863 7046
rect 4887 7044 4943 7046
rect 10229 10906 10285 10908
rect 10309 10906 10365 10908
rect 10389 10906 10445 10908
rect 10469 10906 10525 10908
rect 10229 10854 10275 10906
rect 10275 10854 10285 10906
rect 10309 10854 10339 10906
rect 10339 10854 10351 10906
rect 10351 10854 10365 10906
rect 10389 10854 10403 10906
rect 10403 10854 10415 10906
rect 10415 10854 10445 10906
rect 10469 10854 10479 10906
rect 10479 10854 10525 10906
rect 10229 10852 10285 10854
rect 10309 10852 10365 10854
rect 10389 10852 10445 10854
rect 10469 10852 10525 10854
rect 9569 10362 9625 10364
rect 9649 10362 9705 10364
rect 9729 10362 9785 10364
rect 9809 10362 9865 10364
rect 9569 10310 9615 10362
rect 9615 10310 9625 10362
rect 9649 10310 9679 10362
rect 9679 10310 9691 10362
rect 9691 10310 9705 10362
rect 9729 10310 9743 10362
rect 9743 10310 9755 10362
rect 9755 10310 9785 10362
rect 9809 10310 9819 10362
rect 9819 10310 9865 10362
rect 9569 10308 9625 10310
rect 9649 10308 9705 10310
rect 9729 10308 9785 10310
rect 9809 10308 9865 10310
rect 7108 9274 7164 9276
rect 7188 9274 7244 9276
rect 7268 9274 7324 9276
rect 7348 9274 7404 9276
rect 7108 9222 7154 9274
rect 7154 9222 7164 9274
rect 7188 9222 7218 9274
rect 7218 9222 7230 9274
rect 7230 9222 7244 9274
rect 7268 9222 7282 9274
rect 7282 9222 7294 9274
rect 7294 9222 7324 9274
rect 7348 9222 7358 9274
rect 7358 9222 7404 9274
rect 7108 9220 7164 9222
rect 7188 9220 7244 9222
rect 7268 9220 7324 9222
rect 7348 9220 7404 9222
rect 7768 9818 7824 9820
rect 7848 9818 7904 9820
rect 7928 9818 7984 9820
rect 8008 9818 8064 9820
rect 7768 9766 7814 9818
rect 7814 9766 7824 9818
rect 7848 9766 7878 9818
rect 7878 9766 7890 9818
rect 7890 9766 7904 9818
rect 7928 9766 7942 9818
rect 7942 9766 7954 9818
rect 7954 9766 7984 9818
rect 8008 9766 8018 9818
rect 8018 9766 8064 9818
rect 7768 9764 7824 9766
rect 7848 9764 7904 9766
rect 7928 9764 7984 9766
rect 8008 9764 8064 9766
rect 7768 8730 7824 8732
rect 7848 8730 7904 8732
rect 7928 8730 7984 8732
rect 8008 8730 8064 8732
rect 7768 8678 7814 8730
rect 7814 8678 7824 8730
rect 7848 8678 7878 8730
rect 7878 8678 7890 8730
rect 7890 8678 7904 8730
rect 7928 8678 7942 8730
rect 7942 8678 7954 8730
rect 7954 8678 7984 8730
rect 8008 8678 8018 8730
rect 8018 8678 8064 8730
rect 7768 8676 7824 8678
rect 7848 8676 7904 8678
rect 7928 8676 7984 8678
rect 8008 8676 8064 8678
rect 7108 8186 7164 8188
rect 7188 8186 7244 8188
rect 7268 8186 7324 8188
rect 7348 8186 7404 8188
rect 7108 8134 7154 8186
rect 7154 8134 7164 8186
rect 7188 8134 7218 8186
rect 7218 8134 7230 8186
rect 7230 8134 7244 8186
rect 7268 8134 7282 8186
rect 7282 8134 7294 8186
rect 7294 8134 7324 8186
rect 7348 8134 7358 8186
rect 7358 8134 7404 8186
rect 7108 8132 7164 8134
rect 7188 8132 7244 8134
rect 7268 8132 7324 8134
rect 7348 8132 7404 8134
rect 5170 6976 5226 7032
rect 5998 6840 6054 6896
rect 5307 6554 5363 6556
rect 5387 6554 5443 6556
rect 5467 6554 5523 6556
rect 5547 6554 5603 6556
rect 5307 6502 5353 6554
rect 5353 6502 5363 6554
rect 5387 6502 5417 6554
rect 5417 6502 5429 6554
rect 5429 6502 5443 6554
rect 5467 6502 5481 6554
rect 5481 6502 5493 6554
rect 5493 6502 5523 6554
rect 5547 6502 5557 6554
rect 5557 6502 5603 6554
rect 5307 6500 5363 6502
rect 5387 6500 5443 6502
rect 5467 6500 5523 6502
rect 5547 6500 5603 6502
rect 2846 5466 2902 5468
rect 2926 5466 2982 5468
rect 3006 5466 3062 5468
rect 3086 5466 3142 5468
rect 2846 5414 2892 5466
rect 2892 5414 2902 5466
rect 2926 5414 2956 5466
rect 2956 5414 2968 5466
rect 2968 5414 2982 5466
rect 3006 5414 3020 5466
rect 3020 5414 3032 5466
rect 3032 5414 3062 5466
rect 3086 5414 3096 5466
rect 3096 5414 3142 5466
rect 2846 5412 2902 5414
rect 2926 5412 2982 5414
rect 3006 5412 3062 5414
rect 3086 5412 3142 5414
rect 846 4936 902 4992
rect 2186 4922 2242 4924
rect 2266 4922 2322 4924
rect 2346 4922 2402 4924
rect 2426 4922 2482 4924
rect 2186 4870 2232 4922
rect 2232 4870 2242 4922
rect 2266 4870 2296 4922
rect 2296 4870 2308 4922
rect 2308 4870 2322 4922
rect 2346 4870 2360 4922
rect 2360 4870 2372 4922
rect 2372 4870 2402 4922
rect 2426 4870 2436 4922
rect 2436 4870 2482 4922
rect 2186 4868 2242 4870
rect 2266 4868 2322 4870
rect 2346 4868 2402 4870
rect 2426 4868 2482 4870
rect 4647 6010 4703 6012
rect 4727 6010 4783 6012
rect 4807 6010 4863 6012
rect 4887 6010 4943 6012
rect 4647 5958 4693 6010
rect 4693 5958 4703 6010
rect 4727 5958 4757 6010
rect 4757 5958 4769 6010
rect 4769 5958 4783 6010
rect 4807 5958 4821 6010
rect 4821 5958 4833 6010
rect 4833 5958 4863 6010
rect 4887 5958 4897 6010
rect 4897 5958 4943 6010
rect 4647 5956 4703 5958
rect 4727 5956 4783 5958
rect 4807 5956 4863 5958
rect 4887 5956 4943 5958
rect 5307 5466 5363 5468
rect 5387 5466 5443 5468
rect 5467 5466 5523 5468
rect 5547 5466 5603 5468
rect 5307 5414 5353 5466
rect 5353 5414 5363 5466
rect 5387 5414 5417 5466
rect 5417 5414 5429 5466
rect 5429 5414 5443 5466
rect 5467 5414 5481 5466
rect 5481 5414 5493 5466
rect 5493 5414 5523 5466
rect 5547 5414 5557 5466
rect 5557 5414 5603 5466
rect 5307 5412 5363 5414
rect 5387 5412 5443 5414
rect 5467 5412 5523 5414
rect 5547 5412 5603 5414
rect 4647 4922 4703 4924
rect 4727 4922 4783 4924
rect 4807 4922 4863 4924
rect 4887 4922 4943 4924
rect 4647 4870 4693 4922
rect 4693 4870 4703 4922
rect 4727 4870 4757 4922
rect 4757 4870 4769 4922
rect 4769 4870 4783 4922
rect 4807 4870 4821 4922
rect 4821 4870 4833 4922
rect 4833 4870 4863 4922
rect 4887 4870 4897 4922
rect 4897 4870 4943 4922
rect 4647 4868 4703 4870
rect 4727 4868 4783 4870
rect 4807 4868 4863 4870
rect 4887 4868 4943 4870
rect 2846 4378 2902 4380
rect 2926 4378 2982 4380
rect 3006 4378 3062 4380
rect 3086 4378 3142 4380
rect 2846 4326 2892 4378
rect 2892 4326 2902 4378
rect 2926 4326 2956 4378
rect 2956 4326 2968 4378
rect 2968 4326 2982 4378
rect 3006 4326 3020 4378
rect 3020 4326 3032 4378
rect 3032 4326 3062 4378
rect 3086 4326 3096 4378
rect 3096 4326 3142 4378
rect 2846 4324 2902 4326
rect 2926 4324 2982 4326
rect 3006 4324 3062 4326
rect 3086 4324 3142 4326
rect 2186 3834 2242 3836
rect 2266 3834 2322 3836
rect 2346 3834 2402 3836
rect 2426 3834 2482 3836
rect 2186 3782 2232 3834
rect 2232 3782 2242 3834
rect 2266 3782 2296 3834
rect 2296 3782 2308 3834
rect 2308 3782 2322 3834
rect 2346 3782 2360 3834
rect 2360 3782 2372 3834
rect 2372 3782 2402 3834
rect 2426 3782 2436 3834
rect 2436 3782 2482 3834
rect 2186 3780 2242 3782
rect 2266 3780 2322 3782
rect 2346 3780 2402 3782
rect 2426 3780 2482 3782
rect 2846 3290 2902 3292
rect 2926 3290 2982 3292
rect 3006 3290 3062 3292
rect 3086 3290 3142 3292
rect 2846 3238 2892 3290
rect 2892 3238 2902 3290
rect 2926 3238 2956 3290
rect 2956 3238 2968 3290
rect 2968 3238 2982 3290
rect 3006 3238 3020 3290
rect 3020 3238 3032 3290
rect 3032 3238 3062 3290
rect 3086 3238 3096 3290
rect 3096 3238 3142 3290
rect 2846 3236 2902 3238
rect 2926 3236 2982 3238
rect 3006 3236 3062 3238
rect 3086 3236 3142 3238
rect 4647 3834 4703 3836
rect 4727 3834 4783 3836
rect 4807 3834 4863 3836
rect 4887 3834 4943 3836
rect 4647 3782 4693 3834
rect 4693 3782 4703 3834
rect 4727 3782 4757 3834
rect 4757 3782 4769 3834
rect 4769 3782 4783 3834
rect 4807 3782 4821 3834
rect 4821 3782 4833 3834
rect 4833 3782 4863 3834
rect 4887 3782 4897 3834
rect 4897 3782 4943 3834
rect 4647 3780 4703 3782
rect 4727 3780 4783 3782
rect 4807 3780 4863 3782
rect 4887 3780 4943 3782
rect 2186 2746 2242 2748
rect 2266 2746 2322 2748
rect 2346 2746 2402 2748
rect 2426 2746 2482 2748
rect 2186 2694 2232 2746
rect 2232 2694 2242 2746
rect 2266 2694 2296 2746
rect 2296 2694 2308 2746
rect 2308 2694 2322 2746
rect 2346 2694 2360 2746
rect 2360 2694 2372 2746
rect 2372 2694 2402 2746
rect 2426 2694 2436 2746
rect 2436 2694 2482 2746
rect 2186 2692 2242 2694
rect 2266 2692 2322 2694
rect 2346 2692 2402 2694
rect 2426 2692 2482 2694
rect 5307 4378 5363 4380
rect 5387 4378 5443 4380
rect 5467 4378 5523 4380
rect 5547 4378 5603 4380
rect 5307 4326 5353 4378
rect 5353 4326 5363 4378
rect 5387 4326 5417 4378
rect 5417 4326 5429 4378
rect 5429 4326 5443 4378
rect 5467 4326 5481 4378
rect 5481 4326 5493 4378
rect 5493 4326 5523 4378
rect 5547 4326 5557 4378
rect 5557 4326 5603 4378
rect 5307 4324 5363 4326
rect 5387 4324 5443 4326
rect 5467 4324 5523 4326
rect 5547 4324 5603 4326
rect 4647 2746 4703 2748
rect 4727 2746 4783 2748
rect 4807 2746 4863 2748
rect 4887 2746 4943 2748
rect 4647 2694 4693 2746
rect 4693 2694 4703 2746
rect 4727 2694 4757 2746
rect 4757 2694 4769 2746
rect 4769 2694 4783 2746
rect 4807 2694 4821 2746
rect 4821 2694 4833 2746
rect 4833 2694 4863 2746
rect 4887 2694 4897 2746
rect 4897 2694 4943 2746
rect 4647 2692 4703 2694
rect 4727 2692 4783 2694
rect 4807 2692 4863 2694
rect 4887 2692 4943 2694
rect 5307 3290 5363 3292
rect 5387 3290 5443 3292
rect 5467 3290 5523 3292
rect 5547 3290 5603 3292
rect 5307 3238 5353 3290
rect 5353 3238 5363 3290
rect 5387 3238 5417 3290
rect 5417 3238 5429 3290
rect 5429 3238 5443 3290
rect 5467 3238 5481 3290
rect 5481 3238 5493 3290
rect 5493 3238 5523 3290
rect 5547 3238 5557 3290
rect 5557 3238 5603 3290
rect 5307 3236 5363 3238
rect 5387 3236 5443 3238
rect 5467 3236 5523 3238
rect 5547 3236 5603 3238
rect 7108 7098 7164 7100
rect 7188 7098 7244 7100
rect 7268 7098 7324 7100
rect 7348 7098 7404 7100
rect 7108 7046 7154 7098
rect 7154 7046 7164 7098
rect 7188 7046 7218 7098
rect 7218 7046 7230 7098
rect 7230 7046 7244 7098
rect 7268 7046 7282 7098
rect 7282 7046 7294 7098
rect 7294 7046 7324 7098
rect 7348 7046 7358 7098
rect 7358 7046 7404 7098
rect 7108 7044 7164 7046
rect 7188 7044 7244 7046
rect 7268 7044 7324 7046
rect 7348 7044 7404 7046
rect 7768 7642 7824 7644
rect 7848 7642 7904 7644
rect 7928 7642 7984 7644
rect 8008 7642 8064 7644
rect 7768 7590 7814 7642
rect 7814 7590 7824 7642
rect 7848 7590 7878 7642
rect 7878 7590 7890 7642
rect 7890 7590 7904 7642
rect 7928 7590 7942 7642
rect 7942 7590 7954 7642
rect 7954 7590 7984 7642
rect 8008 7590 8018 7642
rect 8018 7590 8064 7642
rect 7768 7588 7824 7590
rect 7848 7588 7904 7590
rect 7928 7588 7984 7590
rect 8008 7588 8064 7590
rect 7286 6840 7342 6896
rect 10229 9818 10285 9820
rect 10309 9818 10365 9820
rect 10389 9818 10445 9820
rect 10469 9818 10525 9820
rect 10229 9766 10275 9818
rect 10275 9766 10285 9818
rect 10309 9766 10339 9818
rect 10339 9766 10351 9818
rect 10351 9766 10365 9818
rect 10389 9766 10403 9818
rect 10403 9766 10415 9818
rect 10415 9766 10445 9818
rect 10469 9766 10479 9818
rect 10479 9766 10525 9818
rect 10229 9764 10285 9766
rect 10309 9764 10365 9766
rect 10389 9764 10445 9766
rect 10469 9764 10525 9766
rect 10598 9560 10654 9616
rect 9569 9274 9625 9276
rect 9649 9274 9705 9276
rect 9729 9274 9785 9276
rect 9809 9274 9865 9276
rect 9569 9222 9615 9274
rect 9615 9222 9625 9274
rect 9649 9222 9679 9274
rect 9679 9222 9691 9274
rect 9691 9222 9705 9274
rect 9729 9222 9743 9274
rect 9743 9222 9755 9274
rect 9755 9222 9785 9274
rect 9809 9222 9819 9274
rect 9819 9222 9865 9274
rect 9569 9220 9625 9222
rect 9649 9220 9705 9222
rect 9729 9220 9785 9222
rect 9809 9220 9865 9222
rect 10598 8880 10654 8936
rect 10229 8730 10285 8732
rect 10309 8730 10365 8732
rect 10389 8730 10445 8732
rect 10469 8730 10525 8732
rect 10229 8678 10275 8730
rect 10275 8678 10285 8730
rect 10309 8678 10339 8730
rect 10339 8678 10351 8730
rect 10351 8678 10365 8730
rect 10389 8678 10403 8730
rect 10403 8678 10415 8730
rect 10415 8678 10445 8730
rect 10469 8678 10479 8730
rect 10479 8678 10525 8730
rect 10229 8676 10285 8678
rect 10309 8676 10365 8678
rect 10389 8676 10445 8678
rect 10469 8676 10525 8678
rect 7768 6554 7824 6556
rect 7848 6554 7904 6556
rect 7928 6554 7984 6556
rect 8008 6554 8064 6556
rect 7768 6502 7814 6554
rect 7814 6502 7824 6554
rect 7848 6502 7878 6554
rect 7878 6502 7890 6554
rect 7890 6502 7904 6554
rect 7928 6502 7942 6554
rect 7942 6502 7954 6554
rect 7954 6502 7984 6554
rect 8008 6502 8018 6554
rect 8018 6502 8064 6554
rect 7768 6500 7824 6502
rect 7848 6500 7904 6502
rect 7928 6500 7984 6502
rect 8008 6500 8064 6502
rect 7108 6010 7164 6012
rect 7188 6010 7244 6012
rect 7268 6010 7324 6012
rect 7348 6010 7404 6012
rect 7108 5958 7154 6010
rect 7154 5958 7164 6010
rect 7188 5958 7218 6010
rect 7218 5958 7230 6010
rect 7230 5958 7244 6010
rect 7268 5958 7282 6010
rect 7282 5958 7294 6010
rect 7294 5958 7324 6010
rect 7348 5958 7358 6010
rect 7358 5958 7404 6010
rect 7108 5956 7164 5958
rect 7188 5956 7244 5958
rect 7268 5956 7324 5958
rect 7348 5956 7404 5958
rect 7108 4922 7164 4924
rect 7188 4922 7244 4924
rect 7268 4922 7324 4924
rect 7348 4922 7404 4924
rect 7108 4870 7154 4922
rect 7154 4870 7164 4922
rect 7188 4870 7218 4922
rect 7218 4870 7230 4922
rect 7230 4870 7244 4922
rect 7268 4870 7282 4922
rect 7282 4870 7294 4922
rect 7294 4870 7324 4922
rect 7348 4870 7358 4922
rect 7358 4870 7404 4922
rect 7108 4868 7164 4870
rect 7188 4868 7244 4870
rect 7268 4868 7324 4870
rect 7348 4868 7404 4870
rect 7768 5466 7824 5468
rect 7848 5466 7904 5468
rect 7928 5466 7984 5468
rect 8008 5466 8064 5468
rect 7768 5414 7814 5466
rect 7814 5414 7824 5466
rect 7848 5414 7878 5466
rect 7878 5414 7890 5466
rect 7890 5414 7904 5466
rect 7928 5414 7942 5466
rect 7942 5414 7954 5466
rect 7954 5414 7984 5466
rect 8008 5414 8018 5466
rect 8018 5414 8064 5466
rect 7768 5412 7824 5414
rect 7848 5412 7904 5414
rect 7928 5412 7984 5414
rect 8008 5412 8064 5414
rect 7768 4378 7824 4380
rect 7848 4378 7904 4380
rect 7928 4378 7984 4380
rect 8008 4378 8064 4380
rect 7768 4326 7814 4378
rect 7814 4326 7824 4378
rect 7848 4326 7878 4378
rect 7878 4326 7890 4378
rect 7890 4326 7904 4378
rect 7928 4326 7942 4378
rect 7942 4326 7954 4378
rect 7954 4326 7984 4378
rect 8008 4326 8018 4378
rect 8018 4326 8064 4378
rect 7768 4324 7824 4326
rect 7848 4324 7904 4326
rect 7928 4324 7984 4326
rect 8008 4324 8064 4326
rect 7108 3834 7164 3836
rect 7188 3834 7244 3836
rect 7268 3834 7324 3836
rect 7348 3834 7404 3836
rect 7108 3782 7154 3834
rect 7154 3782 7164 3834
rect 7188 3782 7218 3834
rect 7218 3782 7230 3834
rect 7230 3782 7244 3834
rect 7268 3782 7282 3834
rect 7282 3782 7294 3834
rect 7294 3782 7324 3834
rect 7348 3782 7358 3834
rect 7358 3782 7404 3834
rect 7108 3780 7164 3782
rect 7188 3780 7244 3782
rect 7268 3780 7324 3782
rect 7348 3780 7404 3782
rect 9569 8186 9625 8188
rect 9649 8186 9705 8188
rect 9729 8186 9785 8188
rect 9809 8186 9865 8188
rect 9569 8134 9615 8186
rect 9615 8134 9625 8186
rect 9649 8134 9679 8186
rect 9679 8134 9691 8186
rect 9691 8134 9705 8186
rect 9729 8134 9743 8186
rect 9743 8134 9755 8186
rect 9755 8134 9785 8186
rect 9809 8134 9819 8186
rect 9819 8134 9865 8186
rect 9569 8132 9625 8134
rect 9649 8132 9705 8134
rect 9729 8132 9785 8134
rect 9809 8132 9865 8134
rect 9569 7098 9625 7100
rect 9649 7098 9705 7100
rect 9729 7098 9785 7100
rect 9809 7098 9865 7100
rect 9569 7046 9615 7098
rect 9615 7046 9625 7098
rect 9649 7046 9679 7098
rect 9679 7046 9691 7098
rect 9691 7046 9705 7098
rect 9729 7046 9743 7098
rect 9743 7046 9755 7098
rect 9755 7046 9785 7098
rect 9809 7046 9819 7098
rect 9819 7046 9865 7098
rect 9569 7044 9625 7046
rect 9649 7044 9705 7046
rect 9729 7044 9785 7046
rect 9809 7044 9865 7046
rect 9569 6010 9625 6012
rect 9649 6010 9705 6012
rect 9729 6010 9785 6012
rect 9809 6010 9865 6012
rect 9569 5958 9615 6010
rect 9615 5958 9625 6010
rect 9649 5958 9679 6010
rect 9679 5958 9691 6010
rect 9691 5958 9705 6010
rect 9729 5958 9743 6010
rect 9743 5958 9755 6010
rect 9755 5958 9785 6010
rect 9809 5958 9819 6010
rect 9819 5958 9865 6010
rect 9569 5956 9625 5958
rect 9649 5956 9705 5958
rect 9729 5956 9785 5958
rect 9809 5956 9865 5958
rect 10229 7642 10285 7644
rect 10309 7642 10365 7644
rect 10389 7642 10445 7644
rect 10469 7642 10525 7644
rect 10229 7590 10275 7642
rect 10275 7590 10285 7642
rect 10309 7590 10339 7642
rect 10339 7590 10351 7642
rect 10351 7590 10365 7642
rect 10389 7590 10403 7642
rect 10403 7590 10415 7642
rect 10415 7590 10445 7642
rect 10469 7590 10479 7642
rect 10479 7590 10525 7642
rect 10229 7588 10285 7590
rect 10309 7588 10365 7590
rect 10389 7588 10445 7590
rect 10469 7588 10525 7590
rect 10229 6554 10285 6556
rect 10309 6554 10365 6556
rect 10389 6554 10445 6556
rect 10469 6554 10525 6556
rect 10229 6502 10275 6554
rect 10275 6502 10285 6554
rect 10309 6502 10339 6554
rect 10339 6502 10351 6554
rect 10351 6502 10365 6554
rect 10389 6502 10403 6554
rect 10403 6502 10415 6554
rect 10415 6502 10445 6554
rect 10469 6502 10479 6554
rect 10479 6502 10525 6554
rect 10229 6500 10285 6502
rect 10309 6500 10365 6502
rect 10389 6500 10445 6502
rect 10469 6500 10525 6502
rect 10229 5466 10285 5468
rect 10309 5466 10365 5468
rect 10389 5466 10445 5468
rect 10469 5466 10525 5468
rect 10229 5414 10275 5466
rect 10275 5414 10285 5466
rect 10309 5414 10339 5466
rect 10339 5414 10351 5466
rect 10351 5414 10365 5466
rect 10389 5414 10403 5466
rect 10403 5414 10415 5466
rect 10415 5414 10445 5466
rect 10469 5414 10479 5466
rect 10479 5414 10525 5466
rect 10229 5412 10285 5414
rect 10309 5412 10365 5414
rect 10389 5412 10445 5414
rect 10469 5412 10525 5414
rect 9569 4922 9625 4924
rect 9649 4922 9705 4924
rect 9729 4922 9785 4924
rect 9809 4922 9865 4924
rect 9569 4870 9615 4922
rect 9615 4870 9625 4922
rect 9649 4870 9679 4922
rect 9679 4870 9691 4922
rect 9691 4870 9705 4922
rect 9729 4870 9743 4922
rect 9743 4870 9755 4922
rect 9755 4870 9785 4922
rect 9809 4870 9819 4922
rect 9819 4870 9865 4922
rect 9569 4868 9625 4870
rect 9649 4868 9705 4870
rect 9729 4868 9785 4870
rect 9809 4868 9865 4870
rect 10598 4800 10654 4856
rect 7768 3290 7824 3292
rect 7848 3290 7904 3292
rect 7928 3290 7984 3292
rect 8008 3290 8064 3292
rect 7768 3238 7814 3290
rect 7814 3238 7824 3290
rect 7848 3238 7878 3290
rect 7878 3238 7890 3290
rect 7890 3238 7904 3290
rect 7928 3238 7942 3290
rect 7942 3238 7954 3290
rect 7954 3238 7984 3290
rect 8008 3238 8018 3290
rect 8018 3238 8064 3290
rect 7768 3236 7824 3238
rect 7848 3236 7904 3238
rect 7928 3236 7984 3238
rect 8008 3236 8064 3238
rect 7108 2746 7164 2748
rect 7188 2746 7244 2748
rect 7268 2746 7324 2748
rect 7348 2746 7404 2748
rect 7108 2694 7154 2746
rect 7154 2694 7164 2746
rect 7188 2694 7218 2746
rect 7218 2694 7230 2746
rect 7230 2694 7244 2746
rect 7268 2694 7282 2746
rect 7282 2694 7294 2746
rect 7294 2694 7324 2746
rect 7348 2694 7358 2746
rect 7358 2694 7404 2746
rect 7108 2692 7164 2694
rect 7188 2692 7244 2694
rect 7268 2692 7324 2694
rect 7348 2692 7404 2694
rect 9569 3834 9625 3836
rect 9649 3834 9705 3836
rect 9729 3834 9785 3836
rect 9809 3834 9865 3836
rect 9569 3782 9615 3834
rect 9615 3782 9625 3834
rect 9649 3782 9679 3834
rect 9679 3782 9691 3834
rect 9691 3782 9705 3834
rect 9729 3782 9743 3834
rect 9743 3782 9755 3834
rect 9755 3782 9785 3834
rect 9809 3782 9819 3834
rect 9819 3782 9865 3834
rect 9569 3780 9625 3782
rect 9649 3780 9705 3782
rect 9729 3780 9785 3782
rect 9809 3780 9865 3782
rect 10229 4378 10285 4380
rect 10309 4378 10365 4380
rect 10389 4378 10445 4380
rect 10469 4378 10525 4380
rect 10229 4326 10275 4378
rect 10275 4326 10285 4378
rect 10309 4326 10339 4378
rect 10339 4326 10351 4378
rect 10351 4326 10365 4378
rect 10389 4326 10403 4378
rect 10403 4326 10415 4378
rect 10415 4326 10445 4378
rect 10469 4326 10479 4378
rect 10479 4326 10525 4378
rect 10229 4324 10285 4326
rect 10309 4324 10365 4326
rect 10389 4324 10445 4326
rect 10469 4324 10525 4326
rect 10598 3476 10600 3496
rect 10600 3476 10652 3496
rect 10652 3476 10654 3496
rect 10598 3440 10654 3476
rect 10229 3290 10285 3292
rect 10309 3290 10365 3292
rect 10389 3290 10445 3292
rect 10469 3290 10525 3292
rect 10229 3238 10275 3290
rect 10275 3238 10285 3290
rect 10309 3238 10339 3290
rect 10339 3238 10351 3290
rect 10351 3238 10365 3290
rect 10389 3238 10403 3290
rect 10403 3238 10415 3290
rect 10415 3238 10445 3290
rect 10469 3238 10479 3290
rect 10479 3238 10525 3290
rect 10229 3236 10285 3238
rect 10309 3236 10365 3238
rect 10389 3236 10445 3238
rect 10469 3236 10525 3238
rect 9569 2746 9625 2748
rect 9649 2746 9705 2748
rect 9729 2746 9785 2748
rect 9809 2746 9865 2748
rect 9569 2694 9615 2746
rect 9615 2694 9625 2746
rect 9649 2694 9679 2746
rect 9679 2694 9691 2746
rect 9691 2694 9705 2746
rect 9729 2694 9743 2746
rect 9743 2694 9755 2746
rect 9755 2694 9785 2746
rect 9809 2694 9819 2746
rect 9819 2694 9865 2746
rect 9569 2692 9625 2694
rect 9649 2692 9705 2694
rect 9729 2692 9785 2694
rect 9809 2692 9865 2694
rect 2846 2202 2902 2204
rect 2926 2202 2982 2204
rect 3006 2202 3062 2204
rect 3086 2202 3142 2204
rect 2846 2150 2892 2202
rect 2892 2150 2902 2202
rect 2926 2150 2956 2202
rect 2956 2150 2968 2202
rect 2968 2150 2982 2202
rect 3006 2150 3020 2202
rect 3020 2150 3032 2202
rect 3032 2150 3062 2202
rect 3086 2150 3096 2202
rect 3096 2150 3142 2202
rect 2846 2148 2902 2150
rect 2926 2148 2982 2150
rect 3006 2148 3062 2150
rect 3086 2148 3142 2150
rect 5307 2202 5363 2204
rect 5387 2202 5443 2204
rect 5467 2202 5523 2204
rect 5547 2202 5603 2204
rect 5307 2150 5353 2202
rect 5353 2150 5363 2202
rect 5387 2150 5417 2202
rect 5417 2150 5429 2202
rect 5429 2150 5443 2202
rect 5467 2150 5481 2202
rect 5481 2150 5493 2202
rect 5493 2150 5523 2202
rect 5547 2150 5557 2202
rect 5557 2150 5603 2202
rect 5307 2148 5363 2150
rect 5387 2148 5443 2150
rect 5467 2148 5523 2150
rect 5547 2148 5603 2150
rect 7768 2202 7824 2204
rect 7848 2202 7904 2204
rect 7928 2202 7984 2204
rect 8008 2202 8064 2204
rect 7768 2150 7814 2202
rect 7814 2150 7824 2202
rect 7848 2150 7878 2202
rect 7878 2150 7890 2202
rect 7890 2150 7904 2202
rect 7928 2150 7942 2202
rect 7942 2150 7954 2202
rect 7954 2150 7984 2202
rect 8008 2150 8018 2202
rect 8018 2150 8064 2202
rect 7768 2148 7824 2150
rect 7848 2148 7904 2150
rect 7928 2148 7984 2150
rect 8008 2148 8064 2150
rect 10229 2202 10285 2204
rect 10309 2202 10365 2204
rect 10389 2202 10445 2204
rect 10469 2202 10525 2204
rect 10229 2150 10275 2202
rect 10275 2150 10285 2202
rect 10309 2150 10339 2202
rect 10339 2150 10351 2202
rect 10351 2150 10365 2202
rect 10389 2150 10403 2202
rect 10403 2150 10415 2202
rect 10415 2150 10445 2202
rect 10469 2150 10479 2202
rect 10479 2150 10525 2202
rect 10229 2148 10285 2150
rect 10309 2148 10365 2150
rect 10389 2148 10445 2150
rect 10469 2148 10525 2150
<< metal3 >>
rect 2836 12000 3152 12001
rect 2836 11936 2842 12000
rect 2906 11936 2922 12000
rect 2986 11936 3002 12000
rect 3066 11936 3082 12000
rect 3146 11936 3152 12000
rect 2836 11935 3152 11936
rect 5297 12000 5613 12001
rect 5297 11936 5303 12000
rect 5367 11936 5383 12000
rect 5447 11936 5463 12000
rect 5527 11936 5543 12000
rect 5607 11936 5613 12000
rect 5297 11935 5613 11936
rect 7758 12000 8074 12001
rect 7758 11936 7764 12000
rect 7828 11936 7844 12000
rect 7908 11936 7924 12000
rect 7988 11936 8004 12000
rect 8068 11936 8074 12000
rect 7758 11935 8074 11936
rect 10219 12000 10535 12001
rect 10219 11936 10225 12000
rect 10289 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10465 12000
rect 10529 11936 10535 12000
rect 10219 11935 10535 11936
rect 2176 11456 2492 11457
rect 2176 11392 2182 11456
rect 2246 11392 2262 11456
rect 2326 11392 2342 11456
rect 2406 11392 2422 11456
rect 2486 11392 2492 11456
rect 2176 11391 2492 11392
rect 4637 11456 4953 11457
rect 4637 11392 4643 11456
rect 4707 11392 4723 11456
rect 4787 11392 4803 11456
rect 4867 11392 4883 11456
rect 4947 11392 4953 11456
rect 4637 11391 4953 11392
rect 7098 11456 7414 11457
rect 7098 11392 7104 11456
rect 7168 11392 7184 11456
rect 7248 11392 7264 11456
rect 7328 11392 7344 11456
rect 7408 11392 7414 11456
rect 7098 11391 7414 11392
rect 9559 11456 9875 11457
rect 9559 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9805 11456
rect 9869 11392 9875 11456
rect 9559 11391 9875 11392
rect 2836 10912 3152 10913
rect 2836 10848 2842 10912
rect 2906 10848 2922 10912
rect 2986 10848 3002 10912
rect 3066 10848 3082 10912
rect 3146 10848 3152 10912
rect 2836 10847 3152 10848
rect 5297 10912 5613 10913
rect 5297 10848 5303 10912
rect 5367 10848 5383 10912
rect 5447 10848 5463 10912
rect 5527 10848 5543 10912
rect 5607 10848 5613 10912
rect 5297 10847 5613 10848
rect 7758 10912 8074 10913
rect 7758 10848 7764 10912
rect 7828 10848 7844 10912
rect 7908 10848 7924 10912
rect 7988 10848 8004 10912
rect 8068 10848 8074 10912
rect 7758 10847 8074 10848
rect 10219 10912 10535 10913
rect 10219 10848 10225 10912
rect 10289 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10465 10912
rect 10529 10848 10535 10912
rect 10219 10847 10535 10848
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 2176 10368 2492 10369
rect 2176 10304 2182 10368
rect 2246 10304 2262 10368
rect 2326 10304 2342 10368
rect 2406 10304 2422 10368
rect 2486 10304 2492 10368
rect 2176 10303 2492 10304
rect 4637 10368 4953 10369
rect 4637 10304 4643 10368
rect 4707 10304 4723 10368
rect 4787 10304 4803 10368
rect 4867 10304 4883 10368
rect 4947 10304 4953 10368
rect 4637 10303 4953 10304
rect 7098 10368 7414 10369
rect 7098 10304 7104 10368
rect 7168 10304 7184 10368
rect 7248 10304 7264 10368
rect 7328 10304 7344 10368
rect 7408 10304 7414 10368
rect 7098 10303 7414 10304
rect 9559 10368 9875 10369
rect 9559 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9805 10368
rect 9869 10304 9875 10368
rect 9559 10303 9875 10304
rect 0 10208 800 10238
rect 2836 9824 3152 9825
rect 2836 9760 2842 9824
rect 2906 9760 2922 9824
rect 2986 9760 3002 9824
rect 3066 9760 3082 9824
rect 3146 9760 3152 9824
rect 2836 9759 3152 9760
rect 5297 9824 5613 9825
rect 5297 9760 5303 9824
rect 5367 9760 5383 9824
rect 5447 9760 5463 9824
rect 5527 9760 5543 9824
rect 5607 9760 5613 9824
rect 5297 9759 5613 9760
rect 7758 9824 8074 9825
rect 7758 9760 7764 9824
rect 7828 9760 7844 9824
rect 7908 9760 7924 9824
rect 7988 9760 8004 9824
rect 8068 9760 8074 9824
rect 7758 9759 8074 9760
rect 10219 9824 10535 9825
rect 10219 9760 10225 9824
rect 10289 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10465 9824
rect 10529 9760 10535 9824
rect 10219 9759 10535 9760
rect 0 9618 800 9648
rect 5758 9618 5764 9620
rect 0 9558 5764 9618
rect 0 9528 800 9558
rect 5758 9556 5764 9558
rect 5828 9556 5834 9620
rect 10593 9618 10659 9621
rect 11322 9618 12122 9648
rect 10593 9616 12122 9618
rect 10593 9560 10598 9616
rect 10654 9560 12122 9616
rect 10593 9558 12122 9560
rect 10593 9555 10659 9558
rect 11322 9528 12122 9558
rect 2176 9280 2492 9281
rect 2176 9216 2182 9280
rect 2246 9216 2262 9280
rect 2326 9216 2342 9280
rect 2406 9216 2422 9280
rect 2486 9216 2492 9280
rect 2176 9215 2492 9216
rect 4637 9280 4953 9281
rect 4637 9216 4643 9280
rect 4707 9216 4723 9280
rect 4787 9216 4803 9280
rect 4867 9216 4883 9280
rect 4947 9216 4953 9280
rect 4637 9215 4953 9216
rect 7098 9280 7414 9281
rect 7098 9216 7104 9280
rect 7168 9216 7184 9280
rect 7248 9216 7264 9280
rect 7328 9216 7344 9280
rect 7408 9216 7414 9280
rect 7098 9215 7414 9216
rect 9559 9280 9875 9281
rect 9559 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9805 9280
rect 9869 9216 9875 9280
rect 9559 9215 9875 9216
rect 10593 8938 10659 8941
rect 11322 8938 12122 8968
rect 10593 8936 12122 8938
rect 10593 8880 10598 8936
rect 10654 8880 12122 8936
rect 10593 8878 12122 8880
rect 10593 8875 10659 8878
rect 11322 8848 12122 8878
rect 2836 8736 3152 8737
rect 2836 8672 2842 8736
rect 2906 8672 2922 8736
rect 2986 8672 3002 8736
rect 3066 8672 3082 8736
rect 3146 8672 3152 8736
rect 2836 8671 3152 8672
rect 5297 8736 5613 8737
rect 5297 8672 5303 8736
rect 5367 8672 5383 8736
rect 5447 8672 5463 8736
rect 5527 8672 5543 8736
rect 5607 8672 5613 8736
rect 5297 8671 5613 8672
rect 7758 8736 8074 8737
rect 7758 8672 7764 8736
rect 7828 8672 7844 8736
rect 7908 8672 7924 8736
rect 7988 8672 8004 8736
rect 8068 8672 8074 8736
rect 7758 8671 8074 8672
rect 10219 8736 10535 8737
rect 10219 8672 10225 8736
rect 10289 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10465 8736
rect 10529 8672 10535 8736
rect 10219 8671 10535 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 2176 8192 2492 8193
rect 2176 8128 2182 8192
rect 2246 8128 2262 8192
rect 2326 8128 2342 8192
rect 2406 8128 2422 8192
rect 2486 8128 2492 8192
rect 2176 8127 2492 8128
rect 4637 8192 4953 8193
rect 4637 8128 4643 8192
rect 4707 8128 4723 8192
rect 4787 8128 4803 8192
rect 4867 8128 4883 8192
rect 4947 8128 4953 8192
rect 4637 8127 4953 8128
rect 7098 8192 7414 8193
rect 7098 8128 7104 8192
rect 7168 8128 7184 8192
rect 7248 8128 7264 8192
rect 7328 8128 7344 8192
rect 7408 8128 7414 8192
rect 7098 8127 7414 8128
rect 9559 8192 9875 8193
rect 9559 8128 9565 8192
rect 9629 8128 9645 8192
rect 9709 8128 9725 8192
rect 9789 8128 9805 8192
rect 9869 8128 9875 8192
rect 9559 8127 9875 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 2836 7648 3152 7649
rect 2836 7584 2842 7648
rect 2906 7584 2922 7648
rect 2986 7584 3002 7648
rect 3066 7584 3082 7648
rect 3146 7584 3152 7648
rect 2836 7583 3152 7584
rect 5297 7648 5613 7649
rect 5297 7584 5303 7648
rect 5367 7584 5383 7648
rect 5447 7584 5463 7648
rect 5527 7584 5543 7648
rect 5607 7584 5613 7648
rect 5297 7583 5613 7584
rect 7758 7648 8074 7649
rect 7758 7584 7764 7648
rect 7828 7584 7844 7648
rect 7908 7584 7924 7648
rect 7988 7584 8004 7648
rect 8068 7584 8074 7648
rect 7758 7583 8074 7584
rect 10219 7648 10535 7649
rect 10219 7584 10225 7648
rect 10289 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10465 7648
rect 10529 7584 10535 7648
rect 10219 7583 10535 7584
rect 0 7488 800 7518
rect 2176 7104 2492 7105
rect 2176 7040 2182 7104
rect 2246 7040 2262 7104
rect 2326 7040 2342 7104
rect 2406 7040 2422 7104
rect 2486 7040 2492 7104
rect 2176 7039 2492 7040
rect 4637 7104 4953 7105
rect 4637 7040 4643 7104
rect 4707 7040 4723 7104
rect 4787 7040 4803 7104
rect 4867 7040 4883 7104
rect 4947 7040 4953 7104
rect 4637 7039 4953 7040
rect 7098 7104 7414 7105
rect 7098 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7344 7104
rect 7408 7040 7414 7104
rect 7098 7039 7414 7040
rect 9559 7104 9875 7105
rect 9559 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9805 7104
rect 9869 7040 9875 7104
rect 9559 7039 9875 7040
rect 5165 7034 5231 7037
rect 5165 7032 6930 7034
rect 5165 6976 5170 7032
rect 5226 6976 6930 7032
rect 5165 6974 6930 6976
rect 5165 6971 5231 6974
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 5758 6836 5764 6900
rect 5828 6898 5834 6900
rect 5993 6898 6059 6901
rect 5828 6896 6059 6898
rect 5828 6840 5998 6896
rect 6054 6840 6059 6896
rect 5828 6838 6059 6840
rect 6870 6898 6930 6974
rect 7281 6898 7347 6901
rect 6870 6896 7347 6898
rect 6870 6840 7286 6896
rect 7342 6840 7347 6896
rect 6870 6838 7347 6840
rect 5828 6836 5834 6838
rect 5993 6835 6059 6838
rect 7281 6835 7347 6838
rect 2836 6560 3152 6561
rect 2836 6496 2842 6560
rect 2906 6496 2922 6560
rect 2986 6496 3002 6560
rect 3066 6496 3082 6560
rect 3146 6496 3152 6560
rect 2836 6495 3152 6496
rect 5297 6560 5613 6561
rect 5297 6496 5303 6560
rect 5367 6496 5383 6560
rect 5447 6496 5463 6560
rect 5527 6496 5543 6560
rect 5607 6496 5613 6560
rect 5297 6495 5613 6496
rect 7758 6560 8074 6561
rect 7758 6496 7764 6560
rect 7828 6496 7844 6560
rect 7908 6496 7924 6560
rect 7988 6496 8004 6560
rect 8068 6496 8074 6560
rect 7758 6495 8074 6496
rect 10219 6560 10535 6561
rect 10219 6496 10225 6560
rect 10289 6496 10305 6560
rect 10369 6496 10385 6560
rect 10449 6496 10465 6560
rect 10529 6496 10535 6560
rect 10219 6495 10535 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 0 6128 800 6158
rect 2176 6016 2492 6017
rect 2176 5952 2182 6016
rect 2246 5952 2262 6016
rect 2326 5952 2342 6016
rect 2406 5952 2422 6016
rect 2486 5952 2492 6016
rect 2176 5951 2492 5952
rect 4637 6016 4953 6017
rect 4637 5952 4643 6016
rect 4707 5952 4723 6016
rect 4787 5952 4803 6016
rect 4867 5952 4883 6016
rect 4947 5952 4953 6016
rect 4637 5951 4953 5952
rect 7098 6016 7414 6017
rect 7098 5952 7104 6016
rect 7168 5952 7184 6016
rect 7248 5952 7264 6016
rect 7328 5952 7344 6016
rect 7408 5952 7414 6016
rect 7098 5951 7414 5952
rect 9559 6016 9875 6017
rect 9559 5952 9565 6016
rect 9629 5952 9645 6016
rect 9709 5952 9725 6016
rect 9789 5952 9805 6016
rect 9869 5952 9875 6016
rect 9559 5951 9875 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 2836 5472 3152 5473
rect 2836 5408 2842 5472
rect 2906 5408 2922 5472
rect 2986 5408 3002 5472
rect 3066 5408 3082 5472
rect 3146 5408 3152 5472
rect 2836 5407 3152 5408
rect 5297 5472 5613 5473
rect 5297 5408 5303 5472
rect 5367 5408 5383 5472
rect 5447 5408 5463 5472
rect 5527 5408 5543 5472
rect 5607 5408 5613 5472
rect 5297 5407 5613 5408
rect 7758 5472 8074 5473
rect 7758 5408 7764 5472
rect 7828 5408 7844 5472
rect 7908 5408 7924 5472
rect 7988 5408 8004 5472
rect 8068 5408 8074 5472
rect 7758 5407 8074 5408
rect 10219 5472 10535 5473
rect 10219 5408 10225 5472
rect 10289 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10465 5472
rect 10529 5408 10535 5472
rect 10219 5407 10535 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 2176 4928 2492 4929
rect 2176 4864 2182 4928
rect 2246 4864 2262 4928
rect 2326 4864 2342 4928
rect 2406 4864 2422 4928
rect 2486 4864 2492 4928
rect 2176 4863 2492 4864
rect 4637 4928 4953 4929
rect 4637 4864 4643 4928
rect 4707 4864 4723 4928
rect 4787 4864 4803 4928
rect 4867 4864 4883 4928
rect 4947 4864 4953 4928
rect 4637 4863 4953 4864
rect 7098 4928 7414 4929
rect 7098 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7344 4928
rect 7408 4864 7414 4928
rect 7098 4863 7414 4864
rect 9559 4928 9875 4929
rect 9559 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9805 4928
rect 9869 4864 9875 4928
rect 9559 4863 9875 4864
rect 10593 4858 10659 4861
rect 11322 4858 12122 4888
rect 10593 4856 12122 4858
rect 10593 4800 10598 4856
rect 10654 4800 12122 4856
rect 10593 4798 12122 4800
rect 0 4768 800 4798
rect 10593 4795 10659 4798
rect 11322 4768 12122 4798
rect 2836 4384 3152 4385
rect 2836 4320 2842 4384
rect 2906 4320 2922 4384
rect 2986 4320 3002 4384
rect 3066 4320 3082 4384
rect 3146 4320 3152 4384
rect 2836 4319 3152 4320
rect 5297 4384 5613 4385
rect 5297 4320 5303 4384
rect 5367 4320 5383 4384
rect 5447 4320 5463 4384
rect 5527 4320 5543 4384
rect 5607 4320 5613 4384
rect 5297 4319 5613 4320
rect 7758 4384 8074 4385
rect 7758 4320 7764 4384
rect 7828 4320 7844 4384
rect 7908 4320 7924 4384
rect 7988 4320 8004 4384
rect 8068 4320 8074 4384
rect 7758 4319 8074 4320
rect 10219 4384 10535 4385
rect 10219 4320 10225 4384
rect 10289 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10465 4384
rect 10529 4320 10535 4384
rect 10219 4319 10535 4320
rect 2176 3840 2492 3841
rect 2176 3776 2182 3840
rect 2246 3776 2262 3840
rect 2326 3776 2342 3840
rect 2406 3776 2422 3840
rect 2486 3776 2492 3840
rect 2176 3775 2492 3776
rect 4637 3840 4953 3841
rect 4637 3776 4643 3840
rect 4707 3776 4723 3840
rect 4787 3776 4803 3840
rect 4867 3776 4883 3840
rect 4947 3776 4953 3840
rect 4637 3775 4953 3776
rect 7098 3840 7414 3841
rect 7098 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7344 3840
rect 7408 3776 7414 3840
rect 7098 3775 7414 3776
rect 9559 3840 9875 3841
rect 9559 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9805 3840
rect 9869 3776 9875 3840
rect 9559 3775 9875 3776
rect 10593 3498 10659 3501
rect 11322 3498 12122 3528
rect 10593 3496 12122 3498
rect 10593 3440 10598 3496
rect 10654 3440 12122 3496
rect 10593 3438 12122 3440
rect 10593 3435 10659 3438
rect 11322 3408 12122 3438
rect 2836 3296 3152 3297
rect 2836 3232 2842 3296
rect 2906 3232 2922 3296
rect 2986 3232 3002 3296
rect 3066 3232 3082 3296
rect 3146 3232 3152 3296
rect 2836 3231 3152 3232
rect 5297 3296 5613 3297
rect 5297 3232 5303 3296
rect 5367 3232 5383 3296
rect 5447 3232 5463 3296
rect 5527 3232 5543 3296
rect 5607 3232 5613 3296
rect 5297 3231 5613 3232
rect 7758 3296 8074 3297
rect 7758 3232 7764 3296
rect 7828 3232 7844 3296
rect 7908 3232 7924 3296
rect 7988 3232 8004 3296
rect 8068 3232 8074 3296
rect 7758 3231 8074 3232
rect 10219 3296 10535 3297
rect 10219 3232 10225 3296
rect 10289 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10465 3296
rect 10529 3232 10535 3296
rect 10219 3231 10535 3232
rect 2176 2752 2492 2753
rect 2176 2688 2182 2752
rect 2246 2688 2262 2752
rect 2326 2688 2342 2752
rect 2406 2688 2422 2752
rect 2486 2688 2492 2752
rect 2176 2687 2492 2688
rect 4637 2752 4953 2753
rect 4637 2688 4643 2752
rect 4707 2688 4723 2752
rect 4787 2688 4803 2752
rect 4867 2688 4883 2752
rect 4947 2688 4953 2752
rect 4637 2687 4953 2688
rect 7098 2752 7414 2753
rect 7098 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7344 2752
rect 7408 2688 7414 2752
rect 7098 2687 7414 2688
rect 9559 2752 9875 2753
rect 9559 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9805 2752
rect 9869 2688 9875 2752
rect 9559 2687 9875 2688
rect 2836 2208 3152 2209
rect 2836 2144 2842 2208
rect 2906 2144 2922 2208
rect 2986 2144 3002 2208
rect 3066 2144 3082 2208
rect 3146 2144 3152 2208
rect 2836 2143 3152 2144
rect 5297 2208 5613 2209
rect 5297 2144 5303 2208
rect 5367 2144 5383 2208
rect 5447 2144 5463 2208
rect 5527 2144 5543 2208
rect 5607 2144 5613 2208
rect 5297 2143 5613 2144
rect 7758 2208 8074 2209
rect 7758 2144 7764 2208
rect 7828 2144 7844 2208
rect 7908 2144 7924 2208
rect 7988 2144 8004 2208
rect 8068 2144 8074 2208
rect 7758 2143 8074 2144
rect 10219 2208 10535 2209
rect 10219 2144 10225 2208
rect 10289 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10465 2208
rect 10529 2144 10535 2208
rect 10219 2143 10535 2144
<< via3 >>
rect 2842 11996 2906 12000
rect 2842 11940 2846 11996
rect 2846 11940 2902 11996
rect 2902 11940 2906 11996
rect 2842 11936 2906 11940
rect 2922 11996 2986 12000
rect 2922 11940 2926 11996
rect 2926 11940 2982 11996
rect 2982 11940 2986 11996
rect 2922 11936 2986 11940
rect 3002 11996 3066 12000
rect 3002 11940 3006 11996
rect 3006 11940 3062 11996
rect 3062 11940 3066 11996
rect 3002 11936 3066 11940
rect 3082 11996 3146 12000
rect 3082 11940 3086 11996
rect 3086 11940 3142 11996
rect 3142 11940 3146 11996
rect 3082 11936 3146 11940
rect 5303 11996 5367 12000
rect 5303 11940 5307 11996
rect 5307 11940 5363 11996
rect 5363 11940 5367 11996
rect 5303 11936 5367 11940
rect 5383 11996 5447 12000
rect 5383 11940 5387 11996
rect 5387 11940 5443 11996
rect 5443 11940 5447 11996
rect 5383 11936 5447 11940
rect 5463 11996 5527 12000
rect 5463 11940 5467 11996
rect 5467 11940 5523 11996
rect 5523 11940 5527 11996
rect 5463 11936 5527 11940
rect 5543 11996 5607 12000
rect 5543 11940 5547 11996
rect 5547 11940 5603 11996
rect 5603 11940 5607 11996
rect 5543 11936 5607 11940
rect 7764 11996 7828 12000
rect 7764 11940 7768 11996
rect 7768 11940 7824 11996
rect 7824 11940 7828 11996
rect 7764 11936 7828 11940
rect 7844 11996 7908 12000
rect 7844 11940 7848 11996
rect 7848 11940 7904 11996
rect 7904 11940 7908 11996
rect 7844 11936 7908 11940
rect 7924 11996 7988 12000
rect 7924 11940 7928 11996
rect 7928 11940 7984 11996
rect 7984 11940 7988 11996
rect 7924 11936 7988 11940
rect 8004 11996 8068 12000
rect 8004 11940 8008 11996
rect 8008 11940 8064 11996
rect 8064 11940 8068 11996
rect 8004 11936 8068 11940
rect 10225 11996 10289 12000
rect 10225 11940 10229 11996
rect 10229 11940 10285 11996
rect 10285 11940 10289 11996
rect 10225 11936 10289 11940
rect 10305 11996 10369 12000
rect 10305 11940 10309 11996
rect 10309 11940 10365 11996
rect 10365 11940 10369 11996
rect 10305 11936 10369 11940
rect 10385 11996 10449 12000
rect 10385 11940 10389 11996
rect 10389 11940 10445 11996
rect 10445 11940 10449 11996
rect 10385 11936 10449 11940
rect 10465 11996 10529 12000
rect 10465 11940 10469 11996
rect 10469 11940 10525 11996
rect 10525 11940 10529 11996
rect 10465 11936 10529 11940
rect 2182 11452 2246 11456
rect 2182 11396 2186 11452
rect 2186 11396 2242 11452
rect 2242 11396 2246 11452
rect 2182 11392 2246 11396
rect 2262 11452 2326 11456
rect 2262 11396 2266 11452
rect 2266 11396 2322 11452
rect 2322 11396 2326 11452
rect 2262 11392 2326 11396
rect 2342 11452 2406 11456
rect 2342 11396 2346 11452
rect 2346 11396 2402 11452
rect 2402 11396 2406 11452
rect 2342 11392 2406 11396
rect 2422 11452 2486 11456
rect 2422 11396 2426 11452
rect 2426 11396 2482 11452
rect 2482 11396 2486 11452
rect 2422 11392 2486 11396
rect 4643 11452 4707 11456
rect 4643 11396 4647 11452
rect 4647 11396 4703 11452
rect 4703 11396 4707 11452
rect 4643 11392 4707 11396
rect 4723 11452 4787 11456
rect 4723 11396 4727 11452
rect 4727 11396 4783 11452
rect 4783 11396 4787 11452
rect 4723 11392 4787 11396
rect 4803 11452 4867 11456
rect 4803 11396 4807 11452
rect 4807 11396 4863 11452
rect 4863 11396 4867 11452
rect 4803 11392 4867 11396
rect 4883 11452 4947 11456
rect 4883 11396 4887 11452
rect 4887 11396 4943 11452
rect 4943 11396 4947 11452
rect 4883 11392 4947 11396
rect 7104 11452 7168 11456
rect 7104 11396 7108 11452
rect 7108 11396 7164 11452
rect 7164 11396 7168 11452
rect 7104 11392 7168 11396
rect 7184 11452 7248 11456
rect 7184 11396 7188 11452
rect 7188 11396 7244 11452
rect 7244 11396 7248 11452
rect 7184 11392 7248 11396
rect 7264 11452 7328 11456
rect 7264 11396 7268 11452
rect 7268 11396 7324 11452
rect 7324 11396 7328 11452
rect 7264 11392 7328 11396
rect 7344 11452 7408 11456
rect 7344 11396 7348 11452
rect 7348 11396 7404 11452
rect 7404 11396 7408 11452
rect 7344 11392 7408 11396
rect 9565 11452 9629 11456
rect 9565 11396 9569 11452
rect 9569 11396 9625 11452
rect 9625 11396 9629 11452
rect 9565 11392 9629 11396
rect 9645 11452 9709 11456
rect 9645 11396 9649 11452
rect 9649 11396 9705 11452
rect 9705 11396 9709 11452
rect 9645 11392 9709 11396
rect 9725 11452 9789 11456
rect 9725 11396 9729 11452
rect 9729 11396 9785 11452
rect 9785 11396 9789 11452
rect 9725 11392 9789 11396
rect 9805 11452 9869 11456
rect 9805 11396 9809 11452
rect 9809 11396 9865 11452
rect 9865 11396 9869 11452
rect 9805 11392 9869 11396
rect 2842 10908 2906 10912
rect 2842 10852 2846 10908
rect 2846 10852 2902 10908
rect 2902 10852 2906 10908
rect 2842 10848 2906 10852
rect 2922 10908 2986 10912
rect 2922 10852 2926 10908
rect 2926 10852 2982 10908
rect 2982 10852 2986 10908
rect 2922 10848 2986 10852
rect 3002 10908 3066 10912
rect 3002 10852 3006 10908
rect 3006 10852 3062 10908
rect 3062 10852 3066 10908
rect 3002 10848 3066 10852
rect 3082 10908 3146 10912
rect 3082 10852 3086 10908
rect 3086 10852 3142 10908
rect 3142 10852 3146 10908
rect 3082 10848 3146 10852
rect 5303 10908 5367 10912
rect 5303 10852 5307 10908
rect 5307 10852 5363 10908
rect 5363 10852 5367 10908
rect 5303 10848 5367 10852
rect 5383 10908 5447 10912
rect 5383 10852 5387 10908
rect 5387 10852 5443 10908
rect 5443 10852 5447 10908
rect 5383 10848 5447 10852
rect 5463 10908 5527 10912
rect 5463 10852 5467 10908
rect 5467 10852 5523 10908
rect 5523 10852 5527 10908
rect 5463 10848 5527 10852
rect 5543 10908 5607 10912
rect 5543 10852 5547 10908
rect 5547 10852 5603 10908
rect 5603 10852 5607 10908
rect 5543 10848 5607 10852
rect 7764 10908 7828 10912
rect 7764 10852 7768 10908
rect 7768 10852 7824 10908
rect 7824 10852 7828 10908
rect 7764 10848 7828 10852
rect 7844 10908 7908 10912
rect 7844 10852 7848 10908
rect 7848 10852 7904 10908
rect 7904 10852 7908 10908
rect 7844 10848 7908 10852
rect 7924 10908 7988 10912
rect 7924 10852 7928 10908
rect 7928 10852 7984 10908
rect 7984 10852 7988 10908
rect 7924 10848 7988 10852
rect 8004 10908 8068 10912
rect 8004 10852 8008 10908
rect 8008 10852 8064 10908
rect 8064 10852 8068 10908
rect 8004 10848 8068 10852
rect 10225 10908 10289 10912
rect 10225 10852 10229 10908
rect 10229 10852 10285 10908
rect 10285 10852 10289 10908
rect 10225 10848 10289 10852
rect 10305 10908 10369 10912
rect 10305 10852 10309 10908
rect 10309 10852 10365 10908
rect 10365 10852 10369 10908
rect 10305 10848 10369 10852
rect 10385 10908 10449 10912
rect 10385 10852 10389 10908
rect 10389 10852 10445 10908
rect 10445 10852 10449 10908
rect 10385 10848 10449 10852
rect 10465 10908 10529 10912
rect 10465 10852 10469 10908
rect 10469 10852 10525 10908
rect 10525 10852 10529 10908
rect 10465 10848 10529 10852
rect 2182 10364 2246 10368
rect 2182 10308 2186 10364
rect 2186 10308 2242 10364
rect 2242 10308 2246 10364
rect 2182 10304 2246 10308
rect 2262 10364 2326 10368
rect 2262 10308 2266 10364
rect 2266 10308 2322 10364
rect 2322 10308 2326 10364
rect 2262 10304 2326 10308
rect 2342 10364 2406 10368
rect 2342 10308 2346 10364
rect 2346 10308 2402 10364
rect 2402 10308 2406 10364
rect 2342 10304 2406 10308
rect 2422 10364 2486 10368
rect 2422 10308 2426 10364
rect 2426 10308 2482 10364
rect 2482 10308 2486 10364
rect 2422 10304 2486 10308
rect 4643 10364 4707 10368
rect 4643 10308 4647 10364
rect 4647 10308 4703 10364
rect 4703 10308 4707 10364
rect 4643 10304 4707 10308
rect 4723 10364 4787 10368
rect 4723 10308 4727 10364
rect 4727 10308 4783 10364
rect 4783 10308 4787 10364
rect 4723 10304 4787 10308
rect 4803 10364 4867 10368
rect 4803 10308 4807 10364
rect 4807 10308 4863 10364
rect 4863 10308 4867 10364
rect 4803 10304 4867 10308
rect 4883 10364 4947 10368
rect 4883 10308 4887 10364
rect 4887 10308 4943 10364
rect 4943 10308 4947 10364
rect 4883 10304 4947 10308
rect 7104 10364 7168 10368
rect 7104 10308 7108 10364
rect 7108 10308 7164 10364
rect 7164 10308 7168 10364
rect 7104 10304 7168 10308
rect 7184 10364 7248 10368
rect 7184 10308 7188 10364
rect 7188 10308 7244 10364
rect 7244 10308 7248 10364
rect 7184 10304 7248 10308
rect 7264 10364 7328 10368
rect 7264 10308 7268 10364
rect 7268 10308 7324 10364
rect 7324 10308 7328 10364
rect 7264 10304 7328 10308
rect 7344 10364 7408 10368
rect 7344 10308 7348 10364
rect 7348 10308 7404 10364
rect 7404 10308 7408 10364
rect 7344 10304 7408 10308
rect 9565 10364 9629 10368
rect 9565 10308 9569 10364
rect 9569 10308 9625 10364
rect 9625 10308 9629 10364
rect 9565 10304 9629 10308
rect 9645 10364 9709 10368
rect 9645 10308 9649 10364
rect 9649 10308 9705 10364
rect 9705 10308 9709 10364
rect 9645 10304 9709 10308
rect 9725 10364 9789 10368
rect 9725 10308 9729 10364
rect 9729 10308 9785 10364
rect 9785 10308 9789 10364
rect 9725 10304 9789 10308
rect 9805 10364 9869 10368
rect 9805 10308 9809 10364
rect 9809 10308 9865 10364
rect 9865 10308 9869 10364
rect 9805 10304 9869 10308
rect 2842 9820 2906 9824
rect 2842 9764 2846 9820
rect 2846 9764 2902 9820
rect 2902 9764 2906 9820
rect 2842 9760 2906 9764
rect 2922 9820 2986 9824
rect 2922 9764 2926 9820
rect 2926 9764 2982 9820
rect 2982 9764 2986 9820
rect 2922 9760 2986 9764
rect 3002 9820 3066 9824
rect 3002 9764 3006 9820
rect 3006 9764 3062 9820
rect 3062 9764 3066 9820
rect 3002 9760 3066 9764
rect 3082 9820 3146 9824
rect 3082 9764 3086 9820
rect 3086 9764 3142 9820
rect 3142 9764 3146 9820
rect 3082 9760 3146 9764
rect 5303 9820 5367 9824
rect 5303 9764 5307 9820
rect 5307 9764 5363 9820
rect 5363 9764 5367 9820
rect 5303 9760 5367 9764
rect 5383 9820 5447 9824
rect 5383 9764 5387 9820
rect 5387 9764 5443 9820
rect 5443 9764 5447 9820
rect 5383 9760 5447 9764
rect 5463 9820 5527 9824
rect 5463 9764 5467 9820
rect 5467 9764 5523 9820
rect 5523 9764 5527 9820
rect 5463 9760 5527 9764
rect 5543 9820 5607 9824
rect 5543 9764 5547 9820
rect 5547 9764 5603 9820
rect 5603 9764 5607 9820
rect 5543 9760 5607 9764
rect 7764 9820 7828 9824
rect 7764 9764 7768 9820
rect 7768 9764 7824 9820
rect 7824 9764 7828 9820
rect 7764 9760 7828 9764
rect 7844 9820 7908 9824
rect 7844 9764 7848 9820
rect 7848 9764 7904 9820
rect 7904 9764 7908 9820
rect 7844 9760 7908 9764
rect 7924 9820 7988 9824
rect 7924 9764 7928 9820
rect 7928 9764 7984 9820
rect 7984 9764 7988 9820
rect 7924 9760 7988 9764
rect 8004 9820 8068 9824
rect 8004 9764 8008 9820
rect 8008 9764 8064 9820
rect 8064 9764 8068 9820
rect 8004 9760 8068 9764
rect 10225 9820 10289 9824
rect 10225 9764 10229 9820
rect 10229 9764 10285 9820
rect 10285 9764 10289 9820
rect 10225 9760 10289 9764
rect 10305 9820 10369 9824
rect 10305 9764 10309 9820
rect 10309 9764 10365 9820
rect 10365 9764 10369 9820
rect 10305 9760 10369 9764
rect 10385 9820 10449 9824
rect 10385 9764 10389 9820
rect 10389 9764 10445 9820
rect 10445 9764 10449 9820
rect 10385 9760 10449 9764
rect 10465 9820 10529 9824
rect 10465 9764 10469 9820
rect 10469 9764 10525 9820
rect 10525 9764 10529 9820
rect 10465 9760 10529 9764
rect 5764 9556 5828 9620
rect 2182 9276 2246 9280
rect 2182 9220 2186 9276
rect 2186 9220 2242 9276
rect 2242 9220 2246 9276
rect 2182 9216 2246 9220
rect 2262 9276 2326 9280
rect 2262 9220 2266 9276
rect 2266 9220 2322 9276
rect 2322 9220 2326 9276
rect 2262 9216 2326 9220
rect 2342 9276 2406 9280
rect 2342 9220 2346 9276
rect 2346 9220 2402 9276
rect 2402 9220 2406 9276
rect 2342 9216 2406 9220
rect 2422 9276 2486 9280
rect 2422 9220 2426 9276
rect 2426 9220 2482 9276
rect 2482 9220 2486 9276
rect 2422 9216 2486 9220
rect 4643 9276 4707 9280
rect 4643 9220 4647 9276
rect 4647 9220 4703 9276
rect 4703 9220 4707 9276
rect 4643 9216 4707 9220
rect 4723 9276 4787 9280
rect 4723 9220 4727 9276
rect 4727 9220 4783 9276
rect 4783 9220 4787 9276
rect 4723 9216 4787 9220
rect 4803 9276 4867 9280
rect 4803 9220 4807 9276
rect 4807 9220 4863 9276
rect 4863 9220 4867 9276
rect 4803 9216 4867 9220
rect 4883 9276 4947 9280
rect 4883 9220 4887 9276
rect 4887 9220 4943 9276
rect 4943 9220 4947 9276
rect 4883 9216 4947 9220
rect 7104 9276 7168 9280
rect 7104 9220 7108 9276
rect 7108 9220 7164 9276
rect 7164 9220 7168 9276
rect 7104 9216 7168 9220
rect 7184 9276 7248 9280
rect 7184 9220 7188 9276
rect 7188 9220 7244 9276
rect 7244 9220 7248 9276
rect 7184 9216 7248 9220
rect 7264 9276 7328 9280
rect 7264 9220 7268 9276
rect 7268 9220 7324 9276
rect 7324 9220 7328 9276
rect 7264 9216 7328 9220
rect 7344 9276 7408 9280
rect 7344 9220 7348 9276
rect 7348 9220 7404 9276
rect 7404 9220 7408 9276
rect 7344 9216 7408 9220
rect 9565 9276 9629 9280
rect 9565 9220 9569 9276
rect 9569 9220 9625 9276
rect 9625 9220 9629 9276
rect 9565 9216 9629 9220
rect 9645 9276 9709 9280
rect 9645 9220 9649 9276
rect 9649 9220 9705 9276
rect 9705 9220 9709 9276
rect 9645 9216 9709 9220
rect 9725 9276 9789 9280
rect 9725 9220 9729 9276
rect 9729 9220 9785 9276
rect 9785 9220 9789 9276
rect 9725 9216 9789 9220
rect 9805 9276 9869 9280
rect 9805 9220 9809 9276
rect 9809 9220 9865 9276
rect 9865 9220 9869 9276
rect 9805 9216 9869 9220
rect 2842 8732 2906 8736
rect 2842 8676 2846 8732
rect 2846 8676 2902 8732
rect 2902 8676 2906 8732
rect 2842 8672 2906 8676
rect 2922 8732 2986 8736
rect 2922 8676 2926 8732
rect 2926 8676 2982 8732
rect 2982 8676 2986 8732
rect 2922 8672 2986 8676
rect 3002 8732 3066 8736
rect 3002 8676 3006 8732
rect 3006 8676 3062 8732
rect 3062 8676 3066 8732
rect 3002 8672 3066 8676
rect 3082 8732 3146 8736
rect 3082 8676 3086 8732
rect 3086 8676 3142 8732
rect 3142 8676 3146 8732
rect 3082 8672 3146 8676
rect 5303 8732 5367 8736
rect 5303 8676 5307 8732
rect 5307 8676 5363 8732
rect 5363 8676 5367 8732
rect 5303 8672 5367 8676
rect 5383 8732 5447 8736
rect 5383 8676 5387 8732
rect 5387 8676 5443 8732
rect 5443 8676 5447 8732
rect 5383 8672 5447 8676
rect 5463 8732 5527 8736
rect 5463 8676 5467 8732
rect 5467 8676 5523 8732
rect 5523 8676 5527 8732
rect 5463 8672 5527 8676
rect 5543 8732 5607 8736
rect 5543 8676 5547 8732
rect 5547 8676 5603 8732
rect 5603 8676 5607 8732
rect 5543 8672 5607 8676
rect 7764 8732 7828 8736
rect 7764 8676 7768 8732
rect 7768 8676 7824 8732
rect 7824 8676 7828 8732
rect 7764 8672 7828 8676
rect 7844 8732 7908 8736
rect 7844 8676 7848 8732
rect 7848 8676 7904 8732
rect 7904 8676 7908 8732
rect 7844 8672 7908 8676
rect 7924 8732 7988 8736
rect 7924 8676 7928 8732
rect 7928 8676 7984 8732
rect 7984 8676 7988 8732
rect 7924 8672 7988 8676
rect 8004 8732 8068 8736
rect 8004 8676 8008 8732
rect 8008 8676 8064 8732
rect 8064 8676 8068 8732
rect 8004 8672 8068 8676
rect 10225 8732 10289 8736
rect 10225 8676 10229 8732
rect 10229 8676 10285 8732
rect 10285 8676 10289 8732
rect 10225 8672 10289 8676
rect 10305 8732 10369 8736
rect 10305 8676 10309 8732
rect 10309 8676 10365 8732
rect 10365 8676 10369 8732
rect 10305 8672 10369 8676
rect 10385 8732 10449 8736
rect 10385 8676 10389 8732
rect 10389 8676 10445 8732
rect 10445 8676 10449 8732
rect 10385 8672 10449 8676
rect 10465 8732 10529 8736
rect 10465 8676 10469 8732
rect 10469 8676 10525 8732
rect 10525 8676 10529 8732
rect 10465 8672 10529 8676
rect 2182 8188 2246 8192
rect 2182 8132 2186 8188
rect 2186 8132 2242 8188
rect 2242 8132 2246 8188
rect 2182 8128 2246 8132
rect 2262 8188 2326 8192
rect 2262 8132 2266 8188
rect 2266 8132 2322 8188
rect 2322 8132 2326 8188
rect 2262 8128 2326 8132
rect 2342 8188 2406 8192
rect 2342 8132 2346 8188
rect 2346 8132 2402 8188
rect 2402 8132 2406 8188
rect 2342 8128 2406 8132
rect 2422 8188 2486 8192
rect 2422 8132 2426 8188
rect 2426 8132 2482 8188
rect 2482 8132 2486 8188
rect 2422 8128 2486 8132
rect 4643 8188 4707 8192
rect 4643 8132 4647 8188
rect 4647 8132 4703 8188
rect 4703 8132 4707 8188
rect 4643 8128 4707 8132
rect 4723 8188 4787 8192
rect 4723 8132 4727 8188
rect 4727 8132 4783 8188
rect 4783 8132 4787 8188
rect 4723 8128 4787 8132
rect 4803 8188 4867 8192
rect 4803 8132 4807 8188
rect 4807 8132 4863 8188
rect 4863 8132 4867 8188
rect 4803 8128 4867 8132
rect 4883 8188 4947 8192
rect 4883 8132 4887 8188
rect 4887 8132 4943 8188
rect 4943 8132 4947 8188
rect 4883 8128 4947 8132
rect 7104 8188 7168 8192
rect 7104 8132 7108 8188
rect 7108 8132 7164 8188
rect 7164 8132 7168 8188
rect 7104 8128 7168 8132
rect 7184 8188 7248 8192
rect 7184 8132 7188 8188
rect 7188 8132 7244 8188
rect 7244 8132 7248 8188
rect 7184 8128 7248 8132
rect 7264 8188 7328 8192
rect 7264 8132 7268 8188
rect 7268 8132 7324 8188
rect 7324 8132 7328 8188
rect 7264 8128 7328 8132
rect 7344 8188 7408 8192
rect 7344 8132 7348 8188
rect 7348 8132 7404 8188
rect 7404 8132 7408 8188
rect 7344 8128 7408 8132
rect 9565 8188 9629 8192
rect 9565 8132 9569 8188
rect 9569 8132 9625 8188
rect 9625 8132 9629 8188
rect 9565 8128 9629 8132
rect 9645 8188 9709 8192
rect 9645 8132 9649 8188
rect 9649 8132 9705 8188
rect 9705 8132 9709 8188
rect 9645 8128 9709 8132
rect 9725 8188 9789 8192
rect 9725 8132 9729 8188
rect 9729 8132 9785 8188
rect 9785 8132 9789 8188
rect 9725 8128 9789 8132
rect 9805 8188 9869 8192
rect 9805 8132 9809 8188
rect 9809 8132 9865 8188
rect 9865 8132 9869 8188
rect 9805 8128 9869 8132
rect 2842 7644 2906 7648
rect 2842 7588 2846 7644
rect 2846 7588 2902 7644
rect 2902 7588 2906 7644
rect 2842 7584 2906 7588
rect 2922 7644 2986 7648
rect 2922 7588 2926 7644
rect 2926 7588 2982 7644
rect 2982 7588 2986 7644
rect 2922 7584 2986 7588
rect 3002 7644 3066 7648
rect 3002 7588 3006 7644
rect 3006 7588 3062 7644
rect 3062 7588 3066 7644
rect 3002 7584 3066 7588
rect 3082 7644 3146 7648
rect 3082 7588 3086 7644
rect 3086 7588 3142 7644
rect 3142 7588 3146 7644
rect 3082 7584 3146 7588
rect 5303 7644 5367 7648
rect 5303 7588 5307 7644
rect 5307 7588 5363 7644
rect 5363 7588 5367 7644
rect 5303 7584 5367 7588
rect 5383 7644 5447 7648
rect 5383 7588 5387 7644
rect 5387 7588 5443 7644
rect 5443 7588 5447 7644
rect 5383 7584 5447 7588
rect 5463 7644 5527 7648
rect 5463 7588 5467 7644
rect 5467 7588 5523 7644
rect 5523 7588 5527 7644
rect 5463 7584 5527 7588
rect 5543 7644 5607 7648
rect 5543 7588 5547 7644
rect 5547 7588 5603 7644
rect 5603 7588 5607 7644
rect 5543 7584 5607 7588
rect 7764 7644 7828 7648
rect 7764 7588 7768 7644
rect 7768 7588 7824 7644
rect 7824 7588 7828 7644
rect 7764 7584 7828 7588
rect 7844 7644 7908 7648
rect 7844 7588 7848 7644
rect 7848 7588 7904 7644
rect 7904 7588 7908 7644
rect 7844 7584 7908 7588
rect 7924 7644 7988 7648
rect 7924 7588 7928 7644
rect 7928 7588 7984 7644
rect 7984 7588 7988 7644
rect 7924 7584 7988 7588
rect 8004 7644 8068 7648
rect 8004 7588 8008 7644
rect 8008 7588 8064 7644
rect 8064 7588 8068 7644
rect 8004 7584 8068 7588
rect 10225 7644 10289 7648
rect 10225 7588 10229 7644
rect 10229 7588 10285 7644
rect 10285 7588 10289 7644
rect 10225 7584 10289 7588
rect 10305 7644 10369 7648
rect 10305 7588 10309 7644
rect 10309 7588 10365 7644
rect 10365 7588 10369 7644
rect 10305 7584 10369 7588
rect 10385 7644 10449 7648
rect 10385 7588 10389 7644
rect 10389 7588 10445 7644
rect 10445 7588 10449 7644
rect 10385 7584 10449 7588
rect 10465 7644 10529 7648
rect 10465 7588 10469 7644
rect 10469 7588 10525 7644
rect 10525 7588 10529 7644
rect 10465 7584 10529 7588
rect 2182 7100 2246 7104
rect 2182 7044 2186 7100
rect 2186 7044 2242 7100
rect 2242 7044 2246 7100
rect 2182 7040 2246 7044
rect 2262 7100 2326 7104
rect 2262 7044 2266 7100
rect 2266 7044 2322 7100
rect 2322 7044 2326 7100
rect 2262 7040 2326 7044
rect 2342 7100 2406 7104
rect 2342 7044 2346 7100
rect 2346 7044 2402 7100
rect 2402 7044 2406 7100
rect 2342 7040 2406 7044
rect 2422 7100 2486 7104
rect 2422 7044 2426 7100
rect 2426 7044 2482 7100
rect 2482 7044 2486 7100
rect 2422 7040 2486 7044
rect 4643 7100 4707 7104
rect 4643 7044 4647 7100
rect 4647 7044 4703 7100
rect 4703 7044 4707 7100
rect 4643 7040 4707 7044
rect 4723 7100 4787 7104
rect 4723 7044 4727 7100
rect 4727 7044 4783 7100
rect 4783 7044 4787 7100
rect 4723 7040 4787 7044
rect 4803 7100 4867 7104
rect 4803 7044 4807 7100
rect 4807 7044 4863 7100
rect 4863 7044 4867 7100
rect 4803 7040 4867 7044
rect 4883 7100 4947 7104
rect 4883 7044 4887 7100
rect 4887 7044 4943 7100
rect 4943 7044 4947 7100
rect 4883 7040 4947 7044
rect 7104 7100 7168 7104
rect 7104 7044 7108 7100
rect 7108 7044 7164 7100
rect 7164 7044 7168 7100
rect 7104 7040 7168 7044
rect 7184 7100 7248 7104
rect 7184 7044 7188 7100
rect 7188 7044 7244 7100
rect 7244 7044 7248 7100
rect 7184 7040 7248 7044
rect 7264 7100 7328 7104
rect 7264 7044 7268 7100
rect 7268 7044 7324 7100
rect 7324 7044 7328 7100
rect 7264 7040 7328 7044
rect 7344 7100 7408 7104
rect 7344 7044 7348 7100
rect 7348 7044 7404 7100
rect 7404 7044 7408 7100
rect 7344 7040 7408 7044
rect 9565 7100 9629 7104
rect 9565 7044 9569 7100
rect 9569 7044 9625 7100
rect 9625 7044 9629 7100
rect 9565 7040 9629 7044
rect 9645 7100 9709 7104
rect 9645 7044 9649 7100
rect 9649 7044 9705 7100
rect 9705 7044 9709 7100
rect 9645 7040 9709 7044
rect 9725 7100 9789 7104
rect 9725 7044 9729 7100
rect 9729 7044 9785 7100
rect 9785 7044 9789 7100
rect 9725 7040 9789 7044
rect 9805 7100 9869 7104
rect 9805 7044 9809 7100
rect 9809 7044 9865 7100
rect 9865 7044 9869 7100
rect 9805 7040 9869 7044
rect 5764 6836 5828 6900
rect 2842 6556 2906 6560
rect 2842 6500 2846 6556
rect 2846 6500 2902 6556
rect 2902 6500 2906 6556
rect 2842 6496 2906 6500
rect 2922 6556 2986 6560
rect 2922 6500 2926 6556
rect 2926 6500 2982 6556
rect 2982 6500 2986 6556
rect 2922 6496 2986 6500
rect 3002 6556 3066 6560
rect 3002 6500 3006 6556
rect 3006 6500 3062 6556
rect 3062 6500 3066 6556
rect 3002 6496 3066 6500
rect 3082 6556 3146 6560
rect 3082 6500 3086 6556
rect 3086 6500 3142 6556
rect 3142 6500 3146 6556
rect 3082 6496 3146 6500
rect 5303 6556 5367 6560
rect 5303 6500 5307 6556
rect 5307 6500 5363 6556
rect 5363 6500 5367 6556
rect 5303 6496 5367 6500
rect 5383 6556 5447 6560
rect 5383 6500 5387 6556
rect 5387 6500 5443 6556
rect 5443 6500 5447 6556
rect 5383 6496 5447 6500
rect 5463 6556 5527 6560
rect 5463 6500 5467 6556
rect 5467 6500 5523 6556
rect 5523 6500 5527 6556
rect 5463 6496 5527 6500
rect 5543 6556 5607 6560
rect 5543 6500 5547 6556
rect 5547 6500 5603 6556
rect 5603 6500 5607 6556
rect 5543 6496 5607 6500
rect 7764 6556 7828 6560
rect 7764 6500 7768 6556
rect 7768 6500 7824 6556
rect 7824 6500 7828 6556
rect 7764 6496 7828 6500
rect 7844 6556 7908 6560
rect 7844 6500 7848 6556
rect 7848 6500 7904 6556
rect 7904 6500 7908 6556
rect 7844 6496 7908 6500
rect 7924 6556 7988 6560
rect 7924 6500 7928 6556
rect 7928 6500 7984 6556
rect 7984 6500 7988 6556
rect 7924 6496 7988 6500
rect 8004 6556 8068 6560
rect 8004 6500 8008 6556
rect 8008 6500 8064 6556
rect 8064 6500 8068 6556
rect 8004 6496 8068 6500
rect 10225 6556 10289 6560
rect 10225 6500 10229 6556
rect 10229 6500 10285 6556
rect 10285 6500 10289 6556
rect 10225 6496 10289 6500
rect 10305 6556 10369 6560
rect 10305 6500 10309 6556
rect 10309 6500 10365 6556
rect 10365 6500 10369 6556
rect 10305 6496 10369 6500
rect 10385 6556 10449 6560
rect 10385 6500 10389 6556
rect 10389 6500 10445 6556
rect 10445 6500 10449 6556
rect 10385 6496 10449 6500
rect 10465 6556 10529 6560
rect 10465 6500 10469 6556
rect 10469 6500 10525 6556
rect 10525 6500 10529 6556
rect 10465 6496 10529 6500
rect 2182 6012 2246 6016
rect 2182 5956 2186 6012
rect 2186 5956 2242 6012
rect 2242 5956 2246 6012
rect 2182 5952 2246 5956
rect 2262 6012 2326 6016
rect 2262 5956 2266 6012
rect 2266 5956 2322 6012
rect 2322 5956 2326 6012
rect 2262 5952 2326 5956
rect 2342 6012 2406 6016
rect 2342 5956 2346 6012
rect 2346 5956 2402 6012
rect 2402 5956 2406 6012
rect 2342 5952 2406 5956
rect 2422 6012 2486 6016
rect 2422 5956 2426 6012
rect 2426 5956 2482 6012
rect 2482 5956 2486 6012
rect 2422 5952 2486 5956
rect 4643 6012 4707 6016
rect 4643 5956 4647 6012
rect 4647 5956 4703 6012
rect 4703 5956 4707 6012
rect 4643 5952 4707 5956
rect 4723 6012 4787 6016
rect 4723 5956 4727 6012
rect 4727 5956 4783 6012
rect 4783 5956 4787 6012
rect 4723 5952 4787 5956
rect 4803 6012 4867 6016
rect 4803 5956 4807 6012
rect 4807 5956 4863 6012
rect 4863 5956 4867 6012
rect 4803 5952 4867 5956
rect 4883 6012 4947 6016
rect 4883 5956 4887 6012
rect 4887 5956 4943 6012
rect 4943 5956 4947 6012
rect 4883 5952 4947 5956
rect 7104 6012 7168 6016
rect 7104 5956 7108 6012
rect 7108 5956 7164 6012
rect 7164 5956 7168 6012
rect 7104 5952 7168 5956
rect 7184 6012 7248 6016
rect 7184 5956 7188 6012
rect 7188 5956 7244 6012
rect 7244 5956 7248 6012
rect 7184 5952 7248 5956
rect 7264 6012 7328 6016
rect 7264 5956 7268 6012
rect 7268 5956 7324 6012
rect 7324 5956 7328 6012
rect 7264 5952 7328 5956
rect 7344 6012 7408 6016
rect 7344 5956 7348 6012
rect 7348 5956 7404 6012
rect 7404 5956 7408 6012
rect 7344 5952 7408 5956
rect 9565 6012 9629 6016
rect 9565 5956 9569 6012
rect 9569 5956 9625 6012
rect 9625 5956 9629 6012
rect 9565 5952 9629 5956
rect 9645 6012 9709 6016
rect 9645 5956 9649 6012
rect 9649 5956 9705 6012
rect 9705 5956 9709 6012
rect 9645 5952 9709 5956
rect 9725 6012 9789 6016
rect 9725 5956 9729 6012
rect 9729 5956 9785 6012
rect 9785 5956 9789 6012
rect 9725 5952 9789 5956
rect 9805 6012 9869 6016
rect 9805 5956 9809 6012
rect 9809 5956 9865 6012
rect 9865 5956 9869 6012
rect 9805 5952 9869 5956
rect 2842 5468 2906 5472
rect 2842 5412 2846 5468
rect 2846 5412 2902 5468
rect 2902 5412 2906 5468
rect 2842 5408 2906 5412
rect 2922 5468 2986 5472
rect 2922 5412 2926 5468
rect 2926 5412 2982 5468
rect 2982 5412 2986 5468
rect 2922 5408 2986 5412
rect 3002 5468 3066 5472
rect 3002 5412 3006 5468
rect 3006 5412 3062 5468
rect 3062 5412 3066 5468
rect 3002 5408 3066 5412
rect 3082 5468 3146 5472
rect 3082 5412 3086 5468
rect 3086 5412 3142 5468
rect 3142 5412 3146 5468
rect 3082 5408 3146 5412
rect 5303 5468 5367 5472
rect 5303 5412 5307 5468
rect 5307 5412 5363 5468
rect 5363 5412 5367 5468
rect 5303 5408 5367 5412
rect 5383 5468 5447 5472
rect 5383 5412 5387 5468
rect 5387 5412 5443 5468
rect 5443 5412 5447 5468
rect 5383 5408 5447 5412
rect 5463 5468 5527 5472
rect 5463 5412 5467 5468
rect 5467 5412 5523 5468
rect 5523 5412 5527 5468
rect 5463 5408 5527 5412
rect 5543 5468 5607 5472
rect 5543 5412 5547 5468
rect 5547 5412 5603 5468
rect 5603 5412 5607 5468
rect 5543 5408 5607 5412
rect 7764 5468 7828 5472
rect 7764 5412 7768 5468
rect 7768 5412 7824 5468
rect 7824 5412 7828 5468
rect 7764 5408 7828 5412
rect 7844 5468 7908 5472
rect 7844 5412 7848 5468
rect 7848 5412 7904 5468
rect 7904 5412 7908 5468
rect 7844 5408 7908 5412
rect 7924 5468 7988 5472
rect 7924 5412 7928 5468
rect 7928 5412 7984 5468
rect 7984 5412 7988 5468
rect 7924 5408 7988 5412
rect 8004 5468 8068 5472
rect 8004 5412 8008 5468
rect 8008 5412 8064 5468
rect 8064 5412 8068 5468
rect 8004 5408 8068 5412
rect 10225 5468 10289 5472
rect 10225 5412 10229 5468
rect 10229 5412 10285 5468
rect 10285 5412 10289 5468
rect 10225 5408 10289 5412
rect 10305 5468 10369 5472
rect 10305 5412 10309 5468
rect 10309 5412 10365 5468
rect 10365 5412 10369 5468
rect 10305 5408 10369 5412
rect 10385 5468 10449 5472
rect 10385 5412 10389 5468
rect 10389 5412 10445 5468
rect 10445 5412 10449 5468
rect 10385 5408 10449 5412
rect 10465 5468 10529 5472
rect 10465 5412 10469 5468
rect 10469 5412 10525 5468
rect 10525 5412 10529 5468
rect 10465 5408 10529 5412
rect 2182 4924 2246 4928
rect 2182 4868 2186 4924
rect 2186 4868 2242 4924
rect 2242 4868 2246 4924
rect 2182 4864 2246 4868
rect 2262 4924 2326 4928
rect 2262 4868 2266 4924
rect 2266 4868 2322 4924
rect 2322 4868 2326 4924
rect 2262 4864 2326 4868
rect 2342 4924 2406 4928
rect 2342 4868 2346 4924
rect 2346 4868 2402 4924
rect 2402 4868 2406 4924
rect 2342 4864 2406 4868
rect 2422 4924 2486 4928
rect 2422 4868 2426 4924
rect 2426 4868 2482 4924
rect 2482 4868 2486 4924
rect 2422 4864 2486 4868
rect 4643 4924 4707 4928
rect 4643 4868 4647 4924
rect 4647 4868 4703 4924
rect 4703 4868 4707 4924
rect 4643 4864 4707 4868
rect 4723 4924 4787 4928
rect 4723 4868 4727 4924
rect 4727 4868 4783 4924
rect 4783 4868 4787 4924
rect 4723 4864 4787 4868
rect 4803 4924 4867 4928
rect 4803 4868 4807 4924
rect 4807 4868 4863 4924
rect 4863 4868 4867 4924
rect 4803 4864 4867 4868
rect 4883 4924 4947 4928
rect 4883 4868 4887 4924
rect 4887 4868 4943 4924
rect 4943 4868 4947 4924
rect 4883 4864 4947 4868
rect 7104 4924 7168 4928
rect 7104 4868 7108 4924
rect 7108 4868 7164 4924
rect 7164 4868 7168 4924
rect 7104 4864 7168 4868
rect 7184 4924 7248 4928
rect 7184 4868 7188 4924
rect 7188 4868 7244 4924
rect 7244 4868 7248 4924
rect 7184 4864 7248 4868
rect 7264 4924 7328 4928
rect 7264 4868 7268 4924
rect 7268 4868 7324 4924
rect 7324 4868 7328 4924
rect 7264 4864 7328 4868
rect 7344 4924 7408 4928
rect 7344 4868 7348 4924
rect 7348 4868 7404 4924
rect 7404 4868 7408 4924
rect 7344 4864 7408 4868
rect 9565 4924 9629 4928
rect 9565 4868 9569 4924
rect 9569 4868 9625 4924
rect 9625 4868 9629 4924
rect 9565 4864 9629 4868
rect 9645 4924 9709 4928
rect 9645 4868 9649 4924
rect 9649 4868 9705 4924
rect 9705 4868 9709 4924
rect 9645 4864 9709 4868
rect 9725 4924 9789 4928
rect 9725 4868 9729 4924
rect 9729 4868 9785 4924
rect 9785 4868 9789 4924
rect 9725 4864 9789 4868
rect 9805 4924 9869 4928
rect 9805 4868 9809 4924
rect 9809 4868 9865 4924
rect 9865 4868 9869 4924
rect 9805 4864 9869 4868
rect 2842 4380 2906 4384
rect 2842 4324 2846 4380
rect 2846 4324 2902 4380
rect 2902 4324 2906 4380
rect 2842 4320 2906 4324
rect 2922 4380 2986 4384
rect 2922 4324 2926 4380
rect 2926 4324 2982 4380
rect 2982 4324 2986 4380
rect 2922 4320 2986 4324
rect 3002 4380 3066 4384
rect 3002 4324 3006 4380
rect 3006 4324 3062 4380
rect 3062 4324 3066 4380
rect 3002 4320 3066 4324
rect 3082 4380 3146 4384
rect 3082 4324 3086 4380
rect 3086 4324 3142 4380
rect 3142 4324 3146 4380
rect 3082 4320 3146 4324
rect 5303 4380 5367 4384
rect 5303 4324 5307 4380
rect 5307 4324 5363 4380
rect 5363 4324 5367 4380
rect 5303 4320 5367 4324
rect 5383 4380 5447 4384
rect 5383 4324 5387 4380
rect 5387 4324 5443 4380
rect 5443 4324 5447 4380
rect 5383 4320 5447 4324
rect 5463 4380 5527 4384
rect 5463 4324 5467 4380
rect 5467 4324 5523 4380
rect 5523 4324 5527 4380
rect 5463 4320 5527 4324
rect 5543 4380 5607 4384
rect 5543 4324 5547 4380
rect 5547 4324 5603 4380
rect 5603 4324 5607 4380
rect 5543 4320 5607 4324
rect 7764 4380 7828 4384
rect 7764 4324 7768 4380
rect 7768 4324 7824 4380
rect 7824 4324 7828 4380
rect 7764 4320 7828 4324
rect 7844 4380 7908 4384
rect 7844 4324 7848 4380
rect 7848 4324 7904 4380
rect 7904 4324 7908 4380
rect 7844 4320 7908 4324
rect 7924 4380 7988 4384
rect 7924 4324 7928 4380
rect 7928 4324 7984 4380
rect 7984 4324 7988 4380
rect 7924 4320 7988 4324
rect 8004 4380 8068 4384
rect 8004 4324 8008 4380
rect 8008 4324 8064 4380
rect 8064 4324 8068 4380
rect 8004 4320 8068 4324
rect 10225 4380 10289 4384
rect 10225 4324 10229 4380
rect 10229 4324 10285 4380
rect 10285 4324 10289 4380
rect 10225 4320 10289 4324
rect 10305 4380 10369 4384
rect 10305 4324 10309 4380
rect 10309 4324 10365 4380
rect 10365 4324 10369 4380
rect 10305 4320 10369 4324
rect 10385 4380 10449 4384
rect 10385 4324 10389 4380
rect 10389 4324 10445 4380
rect 10445 4324 10449 4380
rect 10385 4320 10449 4324
rect 10465 4380 10529 4384
rect 10465 4324 10469 4380
rect 10469 4324 10525 4380
rect 10525 4324 10529 4380
rect 10465 4320 10529 4324
rect 2182 3836 2246 3840
rect 2182 3780 2186 3836
rect 2186 3780 2242 3836
rect 2242 3780 2246 3836
rect 2182 3776 2246 3780
rect 2262 3836 2326 3840
rect 2262 3780 2266 3836
rect 2266 3780 2322 3836
rect 2322 3780 2326 3836
rect 2262 3776 2326 3780
rect 2342 3836 2406 3840
rect 2342 3780 2346 3836
rect 2346 3780 2402 3836
rect 2402 3780 2406 3836
rect 2342 3776 2406 3780
rect 2422 3836 2486 3840
rect 2422 3780 2426 3836
rect 2426 3780 2482 3836
rect 2482 3780 2486 3836
rect 2422 3776 2486 3780
rect 4643 3836 4707 3840
rect 4643 3780 4647 3836
rect 4647 3780 4703 3836
rect 4703 3780 4707 3836
rect 4643 3776 4707 3780
rect 4723 3836 4787 3840
rect 4723 3780 4727 3836
rect 4727 3780 4783 3836
rect 4783 3780 4787 3836
rect 4723 3776 4787 3780
rect 4803 3836 4867 3840
rect 4803 3780 4807 3836
rect 4807 3780 4863 3836
rect 4863 3780 4867 3836
rect 4803 3776 4867 3780
rect 4883 3836 4947 3840
rect 4883 3780 4887 3836
rect 4887 3780 4943 3836
rect 4943 3780 4947 3836
rect 4883 3776 4947 3780
rect 7104 3836 7168 3840
rect 7104 3780 7108 3836
rect 7108 3780 7164 3836
rect 7164 3780 7168 3836
rect 7104 3776 7168 3780
rect 7184 3836 7248 3840
rect 7184 3780 7188 3836
rect 7188 3780 7244 3836
rect 7244 3780 7248 3836
rect 7184 3776 7248 3780
rect 7264 3836 7328 3840
rect 7264 3780 7268 3836
rect 7268 3780 7324 3836
rect 7324 3780 7328 3836
rect 7264 3776 7328 3780
rect 7344 3836 7408 3840
rect 7344 3780 7348 3836
rect 7348 3780 7404 3836
rect 7404 3780 7408 3836
rect 7344 3776 7408 3780
rect 9565 3836 9629 3840
rect 9565 3780 9569 3836
rect 9569 3780 9625 3836
rect 9625 3780 9629 3836
rect 9565 3776 9629 3780
rect 9645 3836 9709 3840
rect 9645 3780 9649 3836
rect 9649 3780 9705 3836
rect 9705 3780 9709 3836
rect 9645 3776 9709 3780
rect 9725 3836 9789 3840
rect 9725 3780 9729 3836
rect 9729 3780 9785 3836
rect 9785 3780 9789 3836
rect 9725 3776 9789 3780
rect 9805 3836 9869 3840
rect 9805 3780 9809 3836
rect 9809 3780 9865 3836
rect 9865 3780 9869 3836
rect 9805 3776 9869 3780
rect 2842 3292 2906 3296
rect 2842 3236 2846 3292
rect 2846 3236 2902 3292
rect 2902 3236 2906 3292
rect 2842 3232 2906 3236
rect 2922 3292 2986 3296
rect 2922 3236 2926 3292
rect 2926 3236 2982 3292
rect 2982 3236 2986 3292
rect 2922 3232 2986 3236
rect 3002 3292 3066 3296
rect 3002 3236 3006 3292
rect 3006 3236 3062 3292
rect 3062 3236 3066 3292
rect 3002 3232 3066 3236
rect 3082 3292 3146 3296
rect 3082 3236 3086 3292
rect 3086 3236 3142 3292
rect 3142 3236 3146 3292
rect 3082 3232 3146 3236
rect 5303 3292 5367 3296
rect 5303 3236 5307 3292
rect 5307 3236 5363 3292
rect 5363 3236 5367 3292
rect 5303 3232 5367 3236
rect 5383 3292 5447 3296
rect 5383 3236 5387 3292
rect 5387 3236 5443 3292
rect 5443 3236 5447 3292
rect 5383 3232 5447 3236
rect 5463 3292 5527 3296
rect 5463 3236 5467 3292
rect 5467 3236 5523 3292
rect 5523 3236 5527 3292
rect 5463 3232 5527 3236
rect 5543 3292 5607 3296
rect 5543 3236 5547 3292
rect 5547 3236 5603 3292
rect 5603 3236 5607 3292
rect 5543 3232 5607 3236
rect 7764 3292 7828 3296
rect 7764 3236 7768 3292
rect 7768 3236 7824 3292
rect 7824 3236 7828 3292
rect 7764 3232 7828 3236
rect 7844 3292 7908 3296
rect 7844 3236 7848 3292
rect 7848 3236 7904 3292
rect 7904 3236 7908 3292
rect 7844 3232 7908 3236
rect 7924 3292 7988 3296
rect 7924 3236 7928 3292
rect 7928 3236 7984 3292
rect 7984 3236 7988 3292
rect 7924 3232 7988 3236
rect 8004 3292 8068 3296
rect 8004 3236 8008 3292
rect 8008 3236 8064 3292
rect 8064 3236 8068 3292
rect 8004 3232 8068 3236
rect 10225 3292 10289 3296
rect 10225 3236 10229 3292
rect 10229 3236 10285 3292
rect 10285 3236 10289 3292
rect 10225 3232 10289 3236
rect 10305 3292 10369 3296
rect 10305 3236 10309 3292
rect 10309 3236 10365 3292
rect 10365 3236 10369 3292
rect 10305 3232 10369 3236
rect 10385 3292 10449 3296
rect 10385 3236 10389 3292
rect 10389 3236 10445 3292
rect 10445 3236 10449 3292
rect 10385 3232 10449 3236
rect 10465 3292 10529 3296
rect 10465 3236 10469 3292
rect 10469 3236 10525 3292
rect 10525 3236 10529 3292
rect 10465 3232 10529 3236
rect 2182 2748 2246 2752
rect 2182 2692 2186 2748
rect 2186 2692 2242 2748
rect 2242 2692 2246 2748
rect 2182 2688 2246 2692
rect 2262 2748 2326 2752
rect 2262 2692 2266 2748
rect 2266 2692 2322 2748
rect 2322 2692 2326 2748
rect 2262 2688 2326 2692
rect 2342 2748 2406 2752
rect 2342 2692 2346 2748
rect 2346 2692 2402 2748
rect 2402 2692 2406 2748
rect 2342 2688 2406 2692
rect 2422 2748 2486 2752
rect 2422 2692 2426 2748
rect 2426 2692 2482 2748
rect 2482 2692 2486 2748
rect 2422 2688 2486 2692
rect 4643 2748 4707 2752
rect 4643 2692 4647 2748
rect 4647 2692 4703 2748
rect 4703 2692 4707 2748
rect 4643 2688 4707 2692
rect 4723 2748 4787 2752
rect 4723 2692 4727 2748
rect 4727 2692 4783 2748
rect 4783 2692 4787 2748
rect 4723 2688 4787 2692
rect 4803 2748 4867 2752
rect 4803 2692 4807 2748
rect 4807 2692 4863 2748
rect 4863 2692 4867 2748
rect 4803 2688 4867 2692
rect 4883 2748 4947 2752
rect 4883 2692 4887 2748
rect 4887 2692 4943 2748
rect 4943 2692 4947 2748
rect 4883 2688 4947 2692
rect 7104 2748 7168 2752
rect 7104 2692 7108 2748
rect 7108 2692 7164 2748
rect 7164 2692 7168 2748
rect 7104 2688 7168 2692
rect 7184 2748 7248 2752
rect 7184 2692 7188 2748
rect 7188 2692 7244 2748
rect 7244 2692 7248 2748
rect 7184 2688 7248 2692
rect 7264 2748 7328 2752
rect 7264 2692 7268 2748
rect 7268 2692 7324 2748
rect 7324 2692 7328 2748
rect 7264 2688 7328 2692
rect 7344 2748 7408 2752
rect 7344 2692 7348 2748
rect 7348 2692 7404 2748
rect 7404 2692 7408 2748
rect 7344 2688 7408 2692
rect 9565 2748 9629 2752
rect 9565 2692 9569 2748
rect 9569 2692 9625 2748
rect 9625 2692 9629 2748
rect 9565 2688 9629 2692
rect 9645 2748 9709 2752
rect 9645 2692 9649 2748
rect 9649 2692 9705 2748
rect 9705 2692 9709 2748
rect 9645 2688 9709 2692
rect 9725 2748 9789 2752
rect 9725 2692 9729 2748
rect 9729 2692 9785 2748
rect 9785 2692 9789 2748
rect 9725 2688 9789 2692
rect 9805 2748 9869 2752
rect 9805 2692 9809 2748
rect 9809 2692 9865 2748
rect 9865 2692 9869 2748
rect 9805 2688 9869 2692
rect 2842 2204 2906 2208
rect 2842 2148 2846 2204
rect 2846 2148 2902 2204
rect 2902 2148 2906 2204
rect 2842 2144 2906 2148
rect 2922 2204 2986 2208
rect 2922 2148 2926 2204
rect 2926 2148 2982 2204
rect 2982 2148 2986 2204
rect 2922 2144 2986 2148
rect 3002 2204 3066 2208
rect 3002 2148 3006 2204
rect 3006 2148 3062 2204
rect 3062 2148 3066 2204
rect 3002 2144 3066 2148
rect 3082 2204 3146 2208
rect 3082 2148 3086 2204
rect 3086 2148 3142 2204
rect 3142 2148 3146 2204
rect 3082 2144 3146 2148
rect 5303 2204 5367 2208
rect 5303 2148 5307 2204
rect 5307 2148 5363 2204
rect 5363 2148 5367 2204
rect 5303 2144 5367 2148
rect 5383 2204 5447 2208
rect 5383 2148 5387 2204
rect 5387 2148 5443 2204
rect 5443 2148 5447 2204
rect 5383 2144 5447 2148
rect 5463 2204 5527 2208
rect 5463 2148 5467 2204
rect 5467 2148 5523 2204
rect 5523 2148 5527 2204
rect 5463 2144 5527 2148
rect 5543 2204 5607 2208
rect 5543 2148 5547 2204
rect 5547 2148 5603 2204
rect 5603 2148 5607 2204
rect 5543 2144 5607 2148
rect 7764 2204 7828 2208
rect 7764 2148 7768 2204
rect 7768 2148 7824 2204
rect 7824 2148 7828 2204
rect 7764 2144 7828 2148
rect 7844 2204 7908 2208
rect 7844 2148 7848 2204
rect 7848 2148 7904 2204
rect 7904 2148 7908 2204
rect 7844 2144 7908 2148
rect 7924 2204 7988 2208
rect 7924 2148 7928 2204
rect 7928 2148 7984 2204
rect 7984 2148 7988 2204
rect 7924 2144 7988 2148
rect 8004 2204 8068 2208
rect 8004 2148 8008 2204
rect 8008 2148 8064 2204
rect 8064 2148 8068 2204
rect 8004 2144 8068 2148
rect 10225 2204 10289 2208
rect 10225 2148 10229 2204
rect 10229 2148 10285 2204
rect 10285 2148 10289 2204
rect 10225 2144 10289 2148
rect 10305 2204 10369 2208
rect 10305 2148 10309 2204
rect 10309 2148 10365 2204
rect 10365 2148 10369 2204
rect 10305 2144 10369 2148
rect 10385 2204 10449 2208
rect 10385 2148 10389 2204
rect 10389 2148 10445 2204
rect 10445 2148 10449 2204
rect 10385 2144 10449 2148
rect 10465 2204 10529 2208
rect 10465 2148 10469 2204
rect 10469 2148 10525 2204
rect 10525 2148 10529 2204
rect 10465 2144 10529 2148
<< metal4 >>
rect 2174 11456 2494 12016
rect 2174 11392 2182 11456
rect 2246 11392 2262 11456
rect 2326 11392 2342 11456
rect 2406 11392 2422 11456
rect 2486 11392 2494 11456
rect 2174 10862 2494 11392
rect 2174 10626 2216 10862
rect 2452 10626 2494 10862
rect 2174 10368 2494 10626
rect 2174 10304 2182 10368
rect 2246 10304 2262 10368
rect 2326 10304 2342 10368
rect 2406 10304 2422 10368
rect 2486 10304 2494 10368
rect 2174 9280 2494 10304
rect 2174 9216 2182 9280
rect 2246 9216 2262 9280
rect 2326 9216 2342 9280
rect 2406 9216 2422 9280
rect 2486 9216 2494 9280
rect 2174 8414 2494 9216
rect 2174 8192 2216 8414
rect 2452 8192 2494 8414
rect 2174 8128 2182 8192
rect 2246 8128 2262 8178
rect 2326 8128 2342 8178
rect 2406 8128 2422 8178
rect 2486 8128 2494 8192
rect 2174 7104 2494 8128
rect 2174 7040 2182 7104
rect 2246 7040 2262 7104
rect 2326 7040 2342 7104
rect 2406 7040 2422 7104
rect 2486 7040 2494 7104
rect 2174 6016 2494 7040
rect 2174 5952 2182 6016
rect 2246 5966 2262 6016
rect 2326 5966 2342 6016
rect 2406 5966 2422 6016
rect 2486 5952 2494 6016
rect 2174 5730 2216 5952
rect 2452 5730 2494 5952
rect 2174 4928 2494 5730
rect 2174 4864 2182 4928
rect 2246 4864 2262 4928
rect 2326 4864 2342 4928
rect 2406 4864 2422 4928
rect 2486 4864 2494 4928
rect 2174 3840 2494 4864
rect 2174 3776 2182 3840
rect 2246 3776 2262 3840
rect 2326 3776 2342 3840
rect 2406 3776 2422 3840
rect 2486 3776 2494 3840
rect 2174 3518 2494 3776
rect 2174 3282 2216 3518
rect 2452 3282 2494 3518
rect 2174 2752 2494 3282
rect 2174 2688 2182 2752
rect 2246 2688 2262 2752
rect 2326 2688 2342 2752
rect 2406 2688 2422 2752
rect 2486 2688 2494 2752
rect 2174 2128 2494 2688
rect 2834 12000 3154 12016
rect 2834 11936 2842 12000
rect 2906 11936 2922 12000
rect 2986 11936 3002 12000
rect 3066 11936 3082 12000
rect 3146 11936 3154 12000
rect 2834 11522 3154 11936
rect 2834 11286 2876 11522
rect 3112 11286 3154 11522
rect 2834 10912 3154 11286
rect 2834 10848 2842 10912
rect 2906 10848 2922 10912
rect 2986 10848 3002 10912
rect 3066 10848 3082 10912
rect 3146 10848 3154 10912
rect 2834 9824 3154 10848
rect 2834 9760 2842 9824
rect 2906 9760 2922 9824
rect 2986 9760 3002 9824
rect 3066 9760 3082 9824
rect 3146 9760 3154 9824
rect 2834 9074 3154 9760
rect 2834 8838 2876 9074
rect 3112 8838 3154 9074
rect 2834 8736 3154 8838
rect 2834 8672 2842 8736
rect 2906 8672 2922 8736
rect 2986 8672 3002 8736
rect 3066 8672 3082 8736
rect 3146 8672 3154 8736
rect 2834 7648 3154 8672
rect 2834 7584 2842 7648
rect 2906 7584 2922 7648
rect 2986 7584 3002 7648
rect 3066 7584 3082 7648
rect 3146 7584 3154 7648
rect 2834 6626 3154 7584
rect 2834 6560 2876 6626
rect 3112 6560 3154 6626
rect 2834 6496 2842 6560
rect 3146 6496 3154 6560
rect 2834 6390 2876 6496
rect 3112 6390 3154 6496
rect 2834 5472 3154 6390
rect 2834 5408 2842 5472
rect 2906 5408 2922 5472
rect 2986 5408 3002 5472
rect 3066 5408 3082 5472
rect 3146 5408 3154 5472
rect 2834 4384 3154 5408
rect 2834 4320 2842 4384
rect 2906 4320 2922 4384
rect 2986 4320 3002 4384
rect 3066 4320 3082 4384
rect 3146 4320 3154 4384
rect 2834 4178 3154 4320
rect 2834 3942 2876 4178
rect 3112 3942 3154 4178
rect 2834 3296 3154 3942
rect 2834 3232 2842 3296
rect 2906 3232 2922 3296
rect 2986 3232 3002 3296
rect 3066 3232 3082 3296
rect 3146 3232 3154 3296
rect 2834 2208 3154 3232
rect 2834 2144 2842 2208
rect 2906 2144 2922 2208
rect 2986 2144 3002 2208
rect 3066 2144 3082 2208
rect 3146 2144 3154 2208
rect 2834 2128 3154 2144
rect 4635 11456 4955 12016
rect 4635 11392 4643 11456
rect 4707 11392 4723 11456
rect 4787 11392 4803 11456
rect 4867 11392 4883 11456
rect 4947 11392 4955 11456
rect 4635 10862 4955 11392
rect 4635 10626 4677 10862
rect 4913 10626 4955 10862
rect 4635 10368 4955 10626
rect 4635 10304 4643 10368
rect 4707 10304 4723 10368
rect 4787 10304 4803 10368
rect 4867 10304 4883 10368
rect 4947 10304 4955 10368
rect 4635 9280 4955 10304
rect 4635 9216 4643 9280
rect 4707 9216 4723 9280
rect 4787 9216 4803 9280
rect 4867 9216 4883 9280
rect 4947 9216 4955 9280
rect 4635 8414 4955 9216
rect 4635 8192 4677 8414
rect 4913 8192 4955 8414
rect 4635 8128 4643 8192
rect 4707 8128 4723 8178
rect 4787 8128 4803 8178
rect 4867 8128 4883 8178
rect 4947 8128 4955 8192
rect 4635 7104 4955 8128
rect 4635 7040 4643 7104
rect 4707 7040 4723 7104
rect 4787 7040 4803 7104
rect 4867 7040 4883 7104
rect 4947 7040 4955 7104
rect 4635 6016 4955 7040
rect 4635 5952 4643 6016
rect 4707 5966 4723 6016
rect 4787 5966 4803 6016
rect 4867 5966 4883 6016
rect 4947 5952 4955 6016
rect 4635 5730 4677 5952
rect 4913 5730 4955 5952
rect 4635 4928 4955 5730
rect 4635 4864 4643 4928
rect 4707 4864 4723 4928
rect 4787 4864 4803 4928
rect 4867 4864 4883 4928
rect 4947 4864 4955 4928
rect 4635 3840 4955 4864
rect 4635 3776 4643 3840
rect 4707 3776 4723 3840
rect 4787 3776 4803 3840
rect 4867 3776 4883 3840
rect 4947 3776 4955 3840
rect 4635 3518 4955 3776
rect 4635 3282 4677 3518
rect 4913 3282 4955 3518
rect 4635 2752 4955 3282
rect 4635 2688 4643 2752
rect 4707 2688 4723 2752
rect 4787 2688 4803 2752
rect 4867 2688 4883 2752
rect 4947 2688 4955 2752
rect 4635 2128 4955 2688
rect 5295 12000 5615 12016
rect 5295 11936 5303 12000
rect 5367 11936 5383 12000
rect 5447 11936 5463 12000
rect 5527 11936 5543 12000
rect 5607 11936 5615 12000
rect 5295 11522 5615 11936
rect 5295 11286 5337 11522
rect 5573 11286 5615 11522
rect 5295 10912 5615 11286
rect 5295 10848 5303 10912
rect 5367 10848 5383 10912
rect 5447 10848 5463 10912
rect 5527 10848 5543 10912
rect 5607 10848 5615 10912
rect 5295 9824 5615 10848
rect 5295 9760 5303 9824
rect 5367 9760 5383 9824
rect 5447 9760 5463 9824
rect 5527 9760 5543 9824
rect 5607 9760 5615 9824
rect 5295 9074 5615 9760
rect 7096 11456 7416 12016
rect 7096 11392 7104 11456
rect 7168 11392 7184 11456
rect 7248 11392 7264 11456
rect 7328 11392 7344 11456
rect 7408 11392 7416 11456
rect 7096 10862 7416 11392
rect 7096 10626 7138 10862
rect 7374 10626 7416 10862
rect 7096 10368 7416 10626
rect 7096 10304 7104 10368
rect 7168 10304 7184 10368
rect 7248 10304 7264 10368
rect 7328 10304 7344 10368
rect 7408 10304 7416 10368
rect 5763 9620 5829 9621
rect 5763 9556 5764 9620
rect 5828 9556 5829 9620
rect 5763 9555 5829 9556
rect 5295 8838 5337 9074
rect 5573 8838 5615 9074
rect 5295 8736 5615 8838
rect 5295 8672 5303 8736
rect 5367 8672 5383 8736
rect 5447 8672 5463 8736
rect 5527 8672 5543 8736
rect 5607 8672 5615 8736
rect 5295 7648 5615 8672
rect 5295 7584 5303 7648
rect 5367 7584 5383 7648
rect 5447 7584 5463 7648
rect 5527 7584 5543 7648
rect 5607 7584 5615 7648
rect 5295 6626 5615 7584
rect 5766 6901 5826 9555
rect 7096 9280 7416 10304
rect 7096 9216 7104 9280
rect 7168 9216 7184 9280
rect 7248 9216 7264 9280
rect 7328 9216 7344 9280
rect 7408 9216 7416 9280
rect 7096 8414 7416 9216
rect 7096 8192 7138 8414
rect 7374 8192 7416 8414
rect 7096 8128 7104 8192
rect 7168 8128 7184 8178
rect 7248 8128 7264 8178
rect 7328 8128 7344 8178
rect 7408 8128 7416 8192
rect 7096 7104 7416 8128
rect 7096 7040 7104 7104
rect 7168 7040 7184 7104
rect 7248 7040 7264 7104
rect 7328 7040 7344 7104
rect 7408 7040 7416 7104
rect 5763 6900 5829 6901
rect 5763 6836 5764 6900
rect 5828 6836 5829 6900
rect 5763 6835 5829 6836
rect 5295 6560 5337 6626
rect 5573 6560 5615 6626
rect 5295 6496 5303 6560
rect 5607 6496 5615 6560
rect 5295 6390 5337 6496
rect 5573 6390 5615 6496
rect 5295 5472 5615 6390
rect 5295 5408 5303 5472
rect 5367 5408 5383 5472
rect 5447 5408 5463 5472
rect 5527 5408 5543 5472
rect 5607 5408 5615 5472
rect 5295 4384 5615 5408
rect 5295 4320 5303 4384
rect 5367 4320 5383 4384
rect 5447 4320 5463 4384
rect 5527 4320 5543 4384
rect 5607 4320 5615 4384
rect 5295 4178 5615 4320
rect 5295 3942 5337 4178
rect 5573 3942 5615 4178
rect 5295 3296 5615 3942
rect 5295 3232 5303 3296
rect 5367 3232 5383 3296
rect 5447 3232 5463 3296
rect 5527 3232 5543 3296
rect 5607 3232 5615 3296
rect 5295 2208 5615 3232
rect 5295 2144 5303 2208
rect 5367 2144 5383 2208
rect 5447 2144 5463 2208
rect 5527 2144 5543 2208
rect 5607 2144 5615 2208
rect 5295 2128 5615 2144
rect 7096 6016 7416 7040
rect 7096 5952 7104 6016
rect 7168 5966 7184 6016
rect 7248 5966 7264 6016
rect 7328 5966 7344 6016
rect 7408 5952 7416 6016
rect 7096 5730 7138 5952
rect 7374 5730 7416 5952
rect 7096 4928 7416 5730
rect 7096 4864 7104 4928
rect 7168 4864 7184 4928
rect 7248 4864 7264 4928
rect 7328 4864 7344 4928
rect 7408 4864 7416 4928
rect 7096 3840 7416 4864
rect 7096 3776 7104 3840
rect 7168 3776 7184 3840
rect 7248 3776 7264 3840
rect 7328 3776 7344 3840
rect 7408 3776 7416 3840
rect 7096 3518 7416 3776
rect 7096 3282 7138 3518
rect 7374 3282 7416 3518
rect 7096 2752 7416 3282
rect 7096 2688 7104 2752
rect 7168 2688 7184 2752
rect 7248 2688 7264 2752
rect 7328 2688 7344 2752
rect 7408 2688 7416 2752
rect 7096 2128 7416 2688
rect 7756 12000 8076 12016
rect 7756 11936 7764 12000
rect 7828 11936 7844 12000
rect 7908 11936 7924 12000
rect 7988 11936 8004 12000
rect 8068 11936 8076 12000
rect 7756 11522 8076 11936
rect 7756 11286 7798 11522
rect 8034 11286 8076 11522
rect 7756 10912 8076 11286
rect 7756 10848 7764 10912
rect 7828 10848 7844 10912
rect 7908 10848 7924 10912
rect 7988 10848 8004 10912
rect 8068 10848 8076 10912
rect 7756 9824 8076 10848
rect 7756 9760 7764 9824
rect 7828 9760 7844 9824
rect 7908 9760 7924 9824
rect 7988 9760 8004 9824
rect 8068 9760 8076 9824
rect 7756 9074 8076 9760
rect 7756 8838 7798 9074
rect 8034 8838 8076 9074
rect 7756 8736 8076 8838
rect 7756 8672 7764 8736
rect 7828 8672 7844 8736
rect 7908 8672 7924 8736
rect 7988 8672 8004 8736
rect 8068 8672 8076 8736
rect 7756 7648 8076 8672
rect 7756 7584 7764 7648
rect 7828 7584 7844 7648
rect 7908 7584 7924 7648
rect 7988 7584 8004 7648
rect 8068 7584 8076 7648
rect 7756 6626 8076 7584
rect 7756 6560 7798 6626
rect 8034 6560 8076 6626
rect 7756 6496 7764 6560
rect 8068 6496 8076 6560
rect 7756 6390 7798 6496
rect 8034 6390 8076 6496
rect 7756 5472 8076 6390
rect 7756 5408 7764 5472
rect 7828 5408 7844 5472
rect 7908 5408 7924 5472
rect 7988 5408 8004 5472
rect 8068 5408 8076 5472
rect 7756 4384 8076 5408
rect 7756 4320 7764 4384
rect 7828 4320 7844 4384
rect 7908 4320 7924 4384
rect 7988 4320 8004 4384
rect 8068 4320 8076 4384
rect 7756 4178 8076 4320
rect 7756 3942 7798 4178
rect 8034 3942 8076 4178
rect 7756 3296 8076 3942
rect 7756 3232 7764 3296
rect 7828 3232 7844 3296
rect 7908 3232 7924 3296
rect 7988 3232 8004 3296
rect 8068 3232 8076 3296
rect 7756 2208 8076 3232
rect 7756 2144 7764 2208
rect 7828 2144 7844 2208
rect 7908 2144 7924 2208
rect 7988 2144 8004 2208
rect 8068 2144 8076 2208
rect 7756 2128 8076 2144
rect 9557 11456 9877 12016
rect 9557 11392 9565 11456
rect 9629 11392 9645 11456
rect 9709 11392 9725 11456
rect 9789 11392 9805 11456
rect 9869 11392 9877 11456
rect 9557 10862 9877 11392
rect 9557 10626 9599 10862
rect 9835 10626 9877 10862
rect 9557 10368 9877 10626
rect 9557 10304 9565 10368
rect 9629 10304 9645 10368
rect 9709 10304 9725 10368
rect 9789 10304 9805 10368
rect 9869 10304 9877 10368
rect 9557 9280 9877 10304
rect 9557 9216 9565 9280
rect 9629 9216 9645 9280
rect 9709 9216 9725 9280
rect 9789 9216 9805 9280
rect 9869 9216 9877 9280
rect 9557 8414 9877 9216
rect 9557 8192 9599 8414
rect 9835 8192 9877 8414
rect 9557 8128 9565 8192
rect 9629 8128 9645 8178
rect 9709 8128 9725 8178
rect 9789 8128 9805 8178
rect 9869 8128 9877 8192
rect 9557 7104 9877 8128
rect 9557 7040 9565 7104
rect 9629 7040 9645 7104
rect 9709 7040 9725 7104
rect 9789 7040 9805 7104
rect 9869 7040 9877 7104
rect 9557 6016 9877 7040
rect 9557 5952 9565 6016
rect 9629 5966 9645 6016
rect 9709 5966 9725 6016
rect 9789 5966 9805 6016
rect 9869 5952 9877 6016
rect 9557 5730 9599 5952
rect 9835 5730 9877 5952
rect 9557 4928 9877 5730
rect 9557 4864 9565 4928
rect 9629 4864 9645 4928
rect 9709 4864 9725 4928
rect 9789 4864 9805 4928
rect 9869 4864 9877 4928
rect 9557 3840 9877 4864
rect 9557 3776 9565 3840
rect 9629 3776 9645 3840
rect 9709 3776 9725 3840
rect 9789 3776 9805 3840
rect 9869 3776 9877 3840
rect 9557 3518 9877 3776
rect 9557 3282 9599 3518
rect 9835 3282 9877 3518
rect 9557 2752 9877 3282
rect 9557 2688 9565 2752
rect 9629 2688 9645 2752
rect 9709 2688 9725 2752
rect 9789 2688 9805 2752
rect 9869 2688 9877 2752
rect 9557 2128 9877 2688
rect 10217 12000 10537 12016
rect 10217 11936 10225 12000
rect 10289 11936 10305 12000
rect 10369 11936 10385 12000
rect 10449 11936 10465 12000
rect 10529 11936 10537 12000
rect 10217 11522 10537 11936
rect 10217 11286 10259 11522
rect 10495 11286 10537 11522
rect 10217 10912 10537 11286
rect 10217 10848 10225 10912
rect 10289 10848 10305 10912
rect 10369 10848 10385 10912
rect 10449 10848 10465 10912
rect 10529 10848 10537 10912
rect 10217 9824 10537 10848
rect 10217 9760 10225 9824
rect 10289 9760 10305 9824
rect 10369 9760 10385 9824
rect 10449 9760 10465 9824
rect 10529 9760 10537 9824
rect 10217 9074 10537 9760
rect 10217 8838 10259 9074
rect 10495 8838 10537 9074
rect 10217 8736 10537 8838
rect 10217 8672 10225 8736
rect 10289 8672 10305 8736
rect 10369 8672 10385 8736
rect 10449 8672 10465 8736
rect 10529 8672 10537 8736
rect 10217 7648 10537 8672
rect 10217 7584 10225 7648
rect 10289 7584 10305 7648
rect 10369 7584 10385 7648
rect 10449 7584 10465 7648
rect 10529 7584 10537 7648
rect 10217 6626 10537 7584
rect 10217 6560 10259 6626
rect 10495 6560 10537 6626
rect 10217 6496 10225 6560
rect 10529 6496 10537 6560
rect 10217 6390 10259 6496
rect 10495 6390 10537 6496
rect 10217 5472 10537 6390
rect 10217 5408 10225 5472
rect 10289 5408 10305 5472
rect 10369 5408 10385 5472
rect 10449 5408 10465 5472
rect 10529 5408 10537 5472
rect 10217 4384 10537 5408
rect 10217 4320 10225 4384
rect 10289 4320 10305 4384
rect 10369 4320 10385 4384
rect 10449 4320 10465 4384
rect 10529 4320 10537 4384
rect 10217 4178 10537 4320
rect 10217 3942 10259 4178
rect 10495 3942 10537 4178
rect 10217 3296 10537 3942
rect 10217 3232 10225 3296
rect 10289 3232 10305 3296
rect 10369 3232 10385 3296
rect 10449 3232 10465 3296
rect 10529 3232 10537 3296
rect 10217 2208 10537 3232
rect 10217 2144 10225 2208
rect 10289 2144 10305 2208
rect 10369 2144 10385 2208
rect 10449 2144 10465 2208
rect 10529 2144 10537 2208
rect 10217 2128 10537 2144
<< via4 >>
rect 2216 10626 2452 10862
rect 2216 8192 2452 8414
rect 2216 8178 2246 8192
rect 2246 8178 2262 8192
rect 2262 8178 2326 8192
rect 2326 8178 2342 8192
rect 2342 8178 2406 8192
rect 2406 8178 2422 8192
rect 2422 8178 2452 8192
rect 2216 5952 2246 5966
rect 2246 5952 2262 5966
rect 2262 5952 2326 5966
rect 2326 5952 2342 5966
rect 2342 5952 2406 5966
rect 2406 5952 2422 5966
rect 2422 5952 2452 5966
rect 2216 5730 2452 5952
rect 2216 3282 2452 3518
rect 2876 11286 3112 11522
rect 2876 8838 3112 9074
rect 2876 6560 3112 6626
rect 2876 6496 2906 6560
rect 2906 6496 2922 6560
rect 2922 6496 2986 6560
rect 2986 6496 3002 6560
rect 3002 6496 3066 6560
rect 3066 6496 3082 6560
rect 3082 6496 3112 6560
rect 2876 6390 3112 6496
rect 2876 3942 3112 4178
rect 4677 10626 4913 10862
rect 4677 8192 4913 8414
rect 4677 8178 4707 8192
rect 4707 8178 4723 8192
rect 4723 8178 4787 8192
rect 4787 8178 4803 8192
rect 4803 8178 4867 8192
rect 4867 8178 4883 8192
rect 4883 8178 4913 8192
rect 4677 5952 4707 5966
rect 4707 5952 4723 5966
rect 4723 5952 4787 5966
rect 4787 5952 4803 5966
rect 4803 5952 4867 5966
rect 4867 5952 4883 5966
rect 4883 5952 4913 5966
rect 4677 5730 4913 5952
rect 4677 3282 4913 3518
rect 5337 11286 5573 11522
rect 7138 10626 7374 10862
rect 5337 8838 5573 9074
rect 7138 8192 7374 8414
rect 7138 8178 7168 8192
rect 7168 8178 7184 8192
rect 7184 8178 7248 8192
rect 7248 8178 7264 8192
rect 7264 8178 7328 8192
rect 7328 8178 7344 8192
rect 7344 8178 7374 8192
rect 5337 6560 5573 6626
rect 5337 6496 5367 6560
rect 5367 6496 5383 6560
rect 5383 6496 5447 6560
rect 5447 6496 5463 6560
rect 5463 6496 5527 6560
rect 5527 6496 5543 6560
rect 5543 6496 5573 6560
rect 5337 6390 5573 6496
rect 5337 3942 5573 4178
rect 7138 5952 7168 5966
rect 7168 5952 7184 5966
rect 7184 5952 7248 5966
rect 7248 5952 7264 5966
rect 7264 5952 7328 5966
rect 7328 5952 7344 5966
rect 7344 5952 7374 5966
rect 7138 5730 7374 5952
rect 7138 3282 7374 3518
rect 7798 11286 8034 11522
rect 7798 8838 8034 9074
rect 7798 6560 8034 6626
rect 7798 6496 7828 6560
rect 7828 6496 7844 6560
rect 7844 6496 7908 6560
rect 7908 6496 7924 6560
rect 7924 6496 7988 6560
rect 7988 6496 8004 6560
rect 8004 6496 8034 6560
rect 7798 6390 8034 6496
rect 7798 3942 8034 4178
rect 9599 10626 9835 10862
rect 9599 8192 9835 8414
rect 9599 8178 9629 8192
rect 9629 8178 9645 8192
rect 9645 8178 9709 8192
rect 9709 8178 9725 8192
rect 9725 8178 9789 8192
rect 9789 8178 9805 8192
rect 9805 8178 9835 8192
rect 9599 5952 9629 5966
rect 9629 5952 9645 5966
rect 9645 5952 9709 5966
rect 9709 5952 9725 5966
rect 9725 5952 9789 5966
rect 9789 5952 9805 5966
rect 9805 5952 9835 5966
rect 9599 5730 9835 5952
rect 9599 3282 9835 3518
rect 10259 11286 10495 11522
rect 10259 8838 10495 9074
rect 10259 6560 10495 6626
rect 10259 6496 10289 6560
rect 10289 6496 10305 6560
rect 10305 6496 10369 6560
rect 10369 6496 10385 6560
rect 10385 6496 10449 6560
rect 10449 6496 10465 6560
rect 10465 6496 10495 6560
rect 10259 6390 10495 6496
rect 10259 3942 10495 4178
<< metal5 >>
rect 1056 11522 10996 11564
rect 1056 11286 2876 11522
rect 3112 11286 5337 11522
rect 5573 11286 7798 11522
rect 8034 11286 10259 11522
rect 10495 11286 10996 11522
rect 1056 11244 10996 11286
rect 1056 10862 10996 10904
rect 1056 10626 2216 10862
rect 2452 10626 4677 10862
rect 4913 10626 7138 10862
rect 7374 10626 9599 10862
rect 9835 10626 10996 10862
rect 1056 10584 10996 10626
rect 1056 9074 10996 9116
rect 1056 8838 2876 9074
rect 3112 8838 5337 9074
rect 5573 8838 7798 9074
rect 8034 8838 10259 9074
rect 10495 8838 10996 9074
rect 1056 8796 10996 8838
rect 1056 8414 10996 8456
rect 1056 8178 2216 8414
rect 2452 8178 4677 8414
rect 4913 8178 7138 8414
rect 7374 8178 9599 8414
rect 9835 8178 10996 8414
rect 1056 8136 10996 8178
rect 1056 6626 10996 6668
rect 1056 6390 2876 6626
rect 3112 6390 5337 6626
rect 5573 6390 7798 6626
rect 8034 6390 10259 6626
rect 10495 6390 10996 6626
rect 1056 6348 10996 6390
rect 1056 5966 10996 6008
rect 1056 5730 2216 5966
rect 2452 5730 4677 5966
rect 4913 5730 7138 5966
rect 7374 5730 9599 5966
rect 9835 5730 10996 5966
rect 1056 5688 10996 5730
rect 1056 4178 10996 4220
rect 1056 3942 2876 4178
rect 3112 3942 5337 4178
rect 5573 3942 7798 4178
rect 8034 3942 10259 4178
rect 10495 3942 10996 4178
rect 1056 3900 10996 3942
rect 1056 3518 10996 3560
rect 1056 3282 2216 3518
rect 2452 3282 4677 3518
rect 4913 3282 7138 3518
rect 7374 3282 9599 3518
rect 9835 3282 10996 3518
rect 1056 3240 10996 3282
use sky130_fd_sc_hd__mux2_1  _072_
timestamp 0
transform -1 0 5704 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _073_
timestamp 0
transform 1 0 6992 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_1  _074_
timestamp 0
transform 1 0 7912 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _075_
timestamp 0
transform 1 0 7360 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 0
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _077_
timestamp 0
transform 1 0 7912 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _078_
timestamp 0
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _079_
timestamp 0
transform 1 0 6440 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _080_
timestamp 0
transform -1 0 4324 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _081_
timestamp 0
transform -1 0 3772 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _082_
timestamp 0
transform -1 0 3680 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _083_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _084_
timestamp 0
transform -1 0 3680 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 0
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _086_
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 0
transform 1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _088_
timestamp 0
transform 1 0 2668 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 0
transform -1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 0
transform -1 0 3772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _092_
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 0
transform -1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _094_
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 0
transform -1 0 5152 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _096_
timestamp 0
transform -1 0 7636 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 0
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _098_
timestamp 0
transform -1 0 8740 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 0
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _100_
timestamp 0
transform -1 0 9568 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 0
transform 1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _102_
timestamp 0
transform 1 0 9844 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 0
transform 1 0 8464 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _104_
timestamp 0
transform -1 0 6808 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _106_
timestamp 0
transform 1 0 4416 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 0
transform -1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _108_
timestamp 0
transform 1 0 2116 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 0
transform 1 0 1840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _110_
timestamp 0
transform 1 0 2208 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 0
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _112_
timestamp 0
transform 1 0 2208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 0
transform 1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _114_
timestamp 0
transform 1 0 2300 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 0
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _116_
timestamp 0
transform -1 0 8740 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _117_
timestamp 0
transform 1 0 7636 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _118_
timestamp 0
transform -1 0 8188 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _119_
timestamp 0
transform -1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _120_
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _121_
timestamp 0
transform -1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _122_
timestamp 0
transform 1 0 8280 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _123_
timestamp 0
transform -1 0 7636 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 0
transform -1 0 6992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _125_
timestamp 0
transform -1 0 9844 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 0
transform 1 0 10396 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _127_
timestamp 0
transform 1 0 7176 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 0
transform -1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 0
transform 1 0 7820 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 0
transform 1 0 6532 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _131_
timestamp 0
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 0
transform 1 0 10396 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _133_
timestamp 0
transform -1 0 5152 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 0
transform -1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _135_
timestamp 0
transform -1 0 4876 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 0
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _137_
timestamp 0
transform -1 0 4600 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 0
transform 1 0 5060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _139_
timestamp 0
transform -1 0 4600 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 0
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 0
transform -1 0 6256 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 0
transform -1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 0
transform 1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _144_
timestamp 0
transform -1 0 9292 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _145_
timestamp 0
transform -1 0 10396 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _146_
timestamp 0
transform -1 0 10396 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _147_
timestamp 0
transform -1 0 10396 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _148_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _149_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _150_
timestamp 0
transform -1 0 10396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _151_
timestamp 0
transform 1 0 4232 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _152_
timestamp 0
transform 1 0 3956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _153_
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _154_
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _155_
timestamp 0
transform -1 0 6900 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _156_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _157_
timestamp 0
transform 1 0 9016 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _158_
timestamp 0
transform 1 0 1748 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _159_
timestamp 0
transform 1 0 1748 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _160_
timestamp 0
transform 1 0 2208 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _161_
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _162_
timestamp 0
transform 1 0 4784 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _163_
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _164_
timestamp 0
transform 1 0 6900 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _165_
timestamp 0
transform 1 0 8004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _166_
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _167_
timestamp 0
transform -1 0 8372 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _168_
timestamp 0
transform -1 0 6808 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _169_
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _170_
timestamp 0
transform 1 0 1564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _171_
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _172_
timestamp 0
transform 1 0 1656 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _173_
timestamp 0
transform 1 0 1932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform -1 0 5244 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform 1 0 7820 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_1  clkload0
timestamp 0
transform 1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23
timestamp 0
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_34
timestamp 0
transform 1 0 4232 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_42
timestamp 0
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_48
timestamp 0
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_62
timestamp 0
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77
timestamp 0
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_103
timestamp 0
transform 1 0 10580 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_26
timestamp 0
transform 1 0 3496 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_36
timestamp 0
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 0
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_74
timestamp 0
transform 1 0 7912 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_91
timestamp 0
transform 1 0 9476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_103
timestamp 0
transform 1 0 10580 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_45
timestamp 0
transform 1 0 5244 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 0
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_23
timestamp 0
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_37
timestamp 0
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_103
timestamp 0
transform 1 0 10580 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_14
timestamp 0
transform 1 0 2392 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_24
timestamp 0
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_37
timestamp 0
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_52
timestamp 0
transform 1 0 5888 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_70
timestamp 0
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_6
timestamp 0
transform 1 0 1656 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_34
timestamp 0
transform 1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_40
timestamp 0
transform 1 0 4784 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_60
timestamp 0
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_79
timestamp 0
transform 1 0 8372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_85
timestamp 0
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_18
timestamp 0
transform 1 0 2760 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_35
timestamp 0
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_45
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_62
timestamp 0
transform 1 0 6808 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_101
timestamp 0
transform 1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_6
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_35
timestamp 0
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_52
timestamp 0
transform 1 0 5888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_52
timestamp 0
transform 1 0 5888 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 0
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_21
timestamp 0
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 0
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 0
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_103
timestamp 0
transform 1 0 10580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_22
timestamp 0
transform 1 0 3128 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_32
timestamp 0
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_50
timestamp 0
transform 1 0 5704 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_58
timestamp 0
transform 1 0 6440 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_62
timestamp 0
transform 1 0 6808 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_74
timestamp 0
transform 1 0 7912 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_93
timestamp 0
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_103
timestamp 0
transform 1 0 10580 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_29
timestamp 0
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_65
timestamp 0
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_80
timestamp 0
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_92
timestamp 0
transform 1 0 9568 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_12
timestamp 0
transform 1 0 2208 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_58
timestamp 0
transform 1 0 6440 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_66
timestamp 0
transform 1 0 7176 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_71
timestamp 0
transform 1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 0
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_102
timestamp 0
transform 1 0 10488 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_38
timestamp 0
transform 1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 0
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_71
timestamp 0
transform 1 0 7636 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_11
timestamp 0
transform 1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_22
timestamp 0
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_45
timestamp 0
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_6
timestamp 0
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_25
timestamp 0
transform 1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_89
timestamp 0
transform 1 0 9292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_101
timestamp 0
transform 1 0 10396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_11
timestamp 0
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_57
timestamp 0
transform 1 0 6348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_61
timestamp 0
transform 1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_103
timestamp 0
transform 1 0 10580 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_29
timestamp 0
transform 1 0 3772 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_37
timestamp 0
transform 1 0 4508 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_41
timestamp 0
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_46
timestamp 0
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 0
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_76
timestamp 0
transform 1 0 8096 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_85
timestamp 0
transform 1 0 8924 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_97
timestamp 0
transform 1 0 10028 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_103
timestamp 0
transform 1 0 10580 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 4508 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 10396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 3956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 5888 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform 1 0 3772 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform 1 0 9844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform -1 0 5336 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform -1 0 8464 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 6440 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform -1 0 5796 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform -1 0 6072 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform -1 0 10396 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform 1 0 9844 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 5980 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform -1 0 6256 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 3772 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 0
transform -1 0 3680 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 0
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 0
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 0
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 0
transform -1 0 6164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 0
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 0
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 0
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 0
transform -1 0 10672 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 0
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_18
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_19
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_20
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_21
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_22
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 10948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_23
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_24
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 10948 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_25
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_26
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 10948 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_27
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_28
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 10948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_29
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_30
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 10948 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_31
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_32
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 10948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_33
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 10948 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_34
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 10948 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_35
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_40
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_41
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_43
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_44
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_45
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_46
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_47
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_48
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_49
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_50
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_51
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_52
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_53
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_54
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_55
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_56
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_57
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_58
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_59
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_60
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_62
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_63
timestamp 0
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_64
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_65
timestamp 0
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
<< labels >>
rlabel metal1 s 6026 11968 6026 11968 4 VGND
rlabel metal1 s 6026 11424 6026 11424 4 VPWR
rlabel metal2 s 6210 10880 6210 10880 4 _000_
rlabel metal1 s 3031 5270 3031 5270 4 _001_
rlabel metal2 s 6394 5474 6394 5474 4 _002_
rlabel metal1 s 4646 5338 4646 5338 4 _003_
rlabel metal2 s 1886 6562 1886 6562 4 _004_
rlabel metal2 s 1978 7650 1978 7650 4 _005_
rlabel metal2 s 1978 9350 1978 9350 4 _006_
rlabel metal2 s 2249 10642 2249 10642 4 _007_
rlabel metal1 s 2111 4182 2111 4182 4 _008_
rlabel metal1 s 2330 3434 2330 3434 4 _009_
rlabel metal1 s 3894 3434 3894 3434 4 _010_
rlabel metal2 s 5101 3094 5101 3094 4 _011_
rlabel metal2 s 5745 3434 5745 3434 4 _012_
rlabel metal2 s 7682 3298 7682 3298 4 _013_
rlabel metal1 s 8367 3026 8367 3026 4 _014_
rlabel metal2 s 9614 4386 9614 4386 4 _015_
rlabel metal1 s 8372 4794 8372 4794 4 _016_
rlabel metal2 s 9062 9180 9062 9180 4 _017_
rlabel metal2 s 8974 10710 8974 10710 4 _018_
rlabel metal1 s 8878 9146 8878 9146 4 _019_
rlabel metal1 s 8878 9520 8878 9520 4 _020_
rlabel metal1 s 10273 5610 10273 5610 4 _021_
rlabel metal2 s 6660 6290 6660 6290 4 _022_
rlabel metal2 s 6665 7378 6665 7378 4 _023_
rlabel metal1 s 10442 6664 10442 6664 4 _024_
rlabel metal1 s 4354 7786 4354 7786 4 _025_
rlabel metal1 s 4140 8058 4140 8058 4 _026_
rlabel metal1 s 4043 10710 4043 10710 4 _027_
rlabel metal1 s 4227 10030 4227 10030 4 _028_
rlabel metal1 s 6470 10710 6470 10710 4 _029_
rlabel metal1 s 8960 8942 8960 8942 4 _030_
rlabel metal1 s 6026 4250 6026 4250 4 _031_
rlabel metal1 s 7728 3026 7728 3026 4 _032_
rlabel metal2 s 8602 3706 8602 3706 4 _033_
rlabel metal1 s 9660 4114 9660 4114 4 _034_
rlabel metal2 s 8694 4828 8694 4828 4 _035_
rlabel metal2 s 6762 4998 6762 4998 4 _036_
rlabel metal1 s 4508 5202 4508 5202 4 _037_
rlabel metal1 s 2116 6290 2116 6290 4 _038_
rlabel metal1 s 2208 7378 2208 7378 4 _039_
rlabel metal2 s 2254 8772 2254 8772 4 _040_
rlabel metal1 s 2438 10234 2438 10234 4 _041_
rlabel metal2 s 8234 10608 8234 10608 4 _042_
rlabel metal2 s 8142 10676 8142 10676 4 _043_
rlabel metal1 s 8326 8976 8326 8976 4 _044_
rlabel metal1 s 8326 9486 8326 9486 4 _045_
rlabel metal2 s 6946 9724 6946 9724 4 _046_
rlabel metal1 s 4232 9486 4232 9486 4 _047_
rlabel metal1 s 9982 5338 9982 5338 4 _048_
rlabel metal1 s 6026 6324 6026 6324 4 _049_
rlabel metal1 s 7728 6970 7728 6970 4 _050_
rlabel metal1 s 9200 7514 9200 7514 4 _051_
rlabel metal1 s 5428 6630 5428 6630 4 _052_
rlabel metal1 s 6302 9044 6302 9044 4 _053_
rlabel metal2 s 4554 10540 4554 10540 4 _054_
rlabel metal1 s 5934 11220 5934 11220 4 _055_
rlabel metal1 s 5980 10778 5980 10778 4 _056_
rlabel metal1 s 7038 9486 7038 9486 4 _057_
rlabel metal2 s 7498 9146 7498 9146 4 _058_
rlabel metal1 s 9890 7514 9890 7514 4 _059_
rlabel metal1 s 8142 8432 8142 8432 4 _060_
rlabel metal1 s 7958 8568 7958 8568 4 _061_
rlabel metal2 s 7590 8670 7590 8670 4 _062_
rlabel metal2 s 3726 6596 3726 6596 4 _063_
rlabel metal1 s 3266 9350 3266 9350 4 _064_
rlabel metal1 s 3174 6630 3174 6630 4 _065_
rlabel metal1 s 4600 2958 4600 2958 4 _066_
rlabel metal2 s 4186 5508 4186 5508 4 _067_
rlabel metal1 s 2438 4590 2438 4590 4 _068_
rlabel metal1 s 2346 3162 2346 3162 4 _069_
rlabel metal2 s 3634 3638 3634 3638 4 _070_
rlabel metal1 s 4692 4250 4692 4250 4 _071_
rlabel metal1 s 5658 8466 5658 8466 4 bit_cnt\[0\]
rlabel metal1 s 7682 8296 7682 8296 4 bit_cnt\[1\]
rlabel metal2 s 7314 9690 7314 9690 4 bit_cnt\[2\]
rlabel metal3 s 5911 6868 5911 6868 4 clk
rlabel metal2 s 5198 7191 5198 7191 4 clknet_0_clk
rlabel metal1 s 4324 3502 4324 3502 4 clknet_1_0__leaf_clk
rlabel metal1 s 6762 5814 6762 5814 4 clknet_1_1__leaf_clk
rlabel metal1 s 7774 11730 7774 11730 4 cs
rlabel metal1 s 3818 5100 3818 5100 4 lfsr_inst.lfsr_out\[0\]
rlabel metal2 s 6210 5950 6210 5950 4 lfsr_inst.lfsr_out\[10\]
rlabel metal1 s 6394 6120 6394 6120 4 lfsr_inst.lfsr_out\[11\]
rlabel metal2 s 4094 6460 4094 6460 4 lfsr_inst.lfsr_out\[12\]
rlabel metal2 s 3634 8228 3634 8228 4 lfsr_inst.lfsr_out\[13\]
rlabel metal2 s 3082 9180 3082 9180 4 lfsr_inst.lfsr_out\[14\]
rlabel metal2 s 3358 10948 3358 10948 4 lfsr_inst.lfsr_out\[15\]
rlabel metal1 s 3772 3978 3772 3978 4 lfsr_inst.lfsr_out\[1\]
rlabel metal1 s 3726 3706 3726 3706 4 lfsr_inst.lfsr_out\[2\]
rlabel metal1 s 5520 3706 5520 3706 4 lfsr_inst.lfsr_out\[3\]
rlabel metal1 s 5934 3162 5934 3162 4 lfsr_inst.lfsr_out\[4\]
rlabel metal2 s 7590 3876 7590 3876 4 lfsr_inst.lfsr_out\[5\]
rlabel metal1 s 9522 3604 9522 3604 4 lfsr_inst.lfsr_out\[6\]
rlabel metal1 s 9522 3162 9522 3162 4 lfsr_inst.lfsr_out\[7\]
rlabel metal1 s 10304 4114 10304 4114 4 lfsr_inst.lfsr_out\[8\]
rlabel metal1 s 7176 4658 7176 4658 4 lfsr_inst.lfsr_out\[9\]
rlabel metal1 s 5106 5712 5106 5712 4 lfsr_inst.load_seed
rlabel metal3 s 1050 5508 1050 5508 4 lfsr_seed[0]
rlabel metal2 s 6486 1588 6486 1588 4 lfsr_seed[10]
rlabel metal3 s 0 6128 800 6248 4 lfsr_seed[11]
port 7 nsew
rlabel metal3 s 1050 6868 1050 6868 4 lfsr_seed[12]
rlabel metal3 s 0 7488 800 7608 4 lfsr_seed[13]
port 9 nsew
rlabel metal3 s 1050 8228 1050 8228 4 lfsr_seed[14]
rlabel metal3 s 0 10208 800 10328 4 lfsr_seed[15]
port 11 nsew
rlabel metal3 s 0 4768 800 4888 4 lfsr_seed[1]
port 12 nsew
rlabel metal2 s 3266 1588 3266 1588 4 lfsr_seed[2]
rlabel metal2 s 3910 1588 3910 1588 4 lfsr_seed[3]
rlabel metal2 s 5198 1588 5198 1588 4 lfsr_seed[4]
rlabel metal2 s 5842 1588 5842 1588 4 lfsr_seed[5]
rlabel metal2 s 7130 1588 7130 1588 4 lfsr_seed[6]
rlabel metal2 s 8418 1588 8418 1588 4 lfsr_seed[7]
rlabel metal3 s 10626 3485 10626 3485 4 lfsr_seed[8]
rlabel metal2 s 10626 4709 10626 4709 4 lfsr_seed[9]
rlabel metal1 s 10580 8602 10580 8602 4 miso
rlabel metal1 s 7866 10166 7866 10166 4 net1
rlabel metal1 s 3266 2618 3266 2618 4 net10
rlabel metal2 s 4186 2856 4186 2856 4 net11
rlabel metal1 s 5244 2618 5244 2618 4 net12
rlabel metal2 s 6118 3332 6118 3332 4 net13
rlabel metal1 s 7130 2618 7130 2618 4 net14
rlabel metal2 s 8510 3332 8510 3332 4 net15
rlabel metal2 s 10442 3808 10442 3808 4 net16
rlabel metal1 s 10396 4794 10396 4794 4 net17
rlabel metal2 s 10442 10404 10442 10404 4 net18
rlabel metal1 s 10672 8466 10672 8466 4 net19
rlabel metal1 s 2392 5542 2392 5542 4 net2
rlabel metal2 s 6486 10880 6486 10880 4 net20
rlabel metal1 s 6486 4114 6486 4114 4 net21
rlabel metal1 s 7130 3162 7130 3162 4 net22
rlabel metal2 s 8970 3910 8970 3910 4 net23
rlabel metal1 s 3174 3162 3174 3162 4 net24
rlabel metal1 s 9844 3706 9844 3706 4 net25
rlabel metal2 s 2898 4794 2898 4794 4 net26
rlabel metal1 s 5152 4250 5152 4250 4 net27
rlabel metal2 s 4002 3536 4002 3536 4 net28
rlabel metal2 s 3634 9520 3634 9520 4 net29
rlabel metal1 s 6440 2618 6440 2618 4 net3
rlabel metal1 s 6624 4590 6624 4590 4 net30
rlabel metal1 s 9844 5202 9844 5202 4 net31
rlabel metal1 s 10672 6290 10672 6290 4 net32
rlabel metal1 s 4186 9622 4186 9622 4 net33
rlabel metal1 s 7728 4794 7728 4794 4 net34
rlabel metal1 s 4692 8874 4692 8874 4 net35
rlabel metal2 s 3818 7684 3818 7684 4 net36
rlabel metal1 s 8510 7718 8510 7718 4 net37
rlabel metal1 s 5014 10710 5014 10710 4 net38
rlabel metal1 s 5290 11322 5290 11322 4 net39
rlabel metal1 s 4692 5746 4692 5746 4 net4
rlabel metal1 s 4002 6358 4002 6358 4 net40
rlabel metal1 s 10580 7174 10580 7174 4 net41
rlabel metal1 s 4968 6834 4968 6834 4 net42
rlabel metal1 s 4784 6970 4784 6970 4 net43
rlabel metal1 s 5612 5338 5612 5338 4 net44
rlabel metal1 s 2852 8466 2852 8466 4 net45
rlabel metal1 s 3220 6426 3220 6426 4 net46
rlabel metal1 s 2116 7174 2116 7174 4 net5
rlabel metal2 s 2714 7616 2714 7616 4 net6
rlabel metal1 s 2714 8364 2714 8364 4 net7
rlabel metal1 s 2208 10098 2208 10098 4 net8
rlabel metal1 s 2898 4658 2898 4658 4 net9
rlabel metal2 s 10626 9809 10626 9809 4 sclk
rlabel metal1 s 7728 10778 7728 10778 4 seeded
rlabel metal1 s 8924 5882 8924 5882 4 tx_buffer\[0\]
rlabel metal1 s 8372 6086 8372 6086 4 tx_buffer\[1\]
rlabel metal1 s 8050 7378 8050 7378 4 tx_buffer\[2\]
rlabel metal1 s 8648 6630 8648 6630 4 tx_buffer\[3\]
rlabel metal1 s 5704 8058 5704 8058 4 tx_buffer\[4\]
rlabel metal1 s 5520 8602 5520 8602 4 tx_buffer\[5\]
rlabel metal1 s 5106 10778 5106 10778 4 tx_buffer\[6\]
rlabel metal2 s 5198 10404 5198 10404 4 tx_buffer\[7\]
flabel metal5 s 1056 11244 10996 11564 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8796 10996 9116 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6348 10996 6668 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3900 10996 4220 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 10217 2128 10537 12016 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7756 2128 8076 12016 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5295 2128 5615 12016 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2834 2128 3154 12016 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 10584 10996 10904 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8136 10996 8456 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5688 10996 6008 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3240 10996 3560 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 9557 2128 9877 12016 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7096 2128 7416 12016 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4635 2128 4955 12016 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2174 2128 2494 12016 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal2 s 7746 13466 7802 14266 0 FreeSans 280 90 0 0 cs
port 4 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 lfsr_seed[0]
port 5 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 lfsr_seed[10]
port 6 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 lfsr_seed[11]
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 lfsr_seed[12]
port 8 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 lfsr_seed[13]
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 lfsr_seed[14]
port 10 nsew
flabel metal3 s 400 10268 400 10268 0 FreeSans 600 0 0 0 lfsr_seed[15]
flabel metal3 s 400 4828 400 4828 0 FreeSans 600 0 0 0 lfsr_seed[1]
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 lfsr_seed[2]
port 13 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 lfsr_seed[3]
port 14 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 lfsr_seed[4]
port 15 nsew
flabel metal2 s 5814 0 5870 800 0 FreeSans 280 90 0 0 lfsr_seed[5]
port 16 nsew
flabel metal2 s 7102 0 7158 800 0 FreeSans 280 90 0 0 lfsr_seed[6]
port 17 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 lfsr_seed[7]
port 18 nsew
flabel metal3 s 11322 3408 12122 3528 0 FreeSans 600 0 0 0 lfsr_seed[8]
port 19 nsew
flabel metal3 s 11322 4768 12122 4888 0 FreeSans 600 0 0 0 lfsr_seed[9]
port 20 nsew
flabel metal3 s 11322 8848 12122 8968 0 FreeSans 600 0 0 0 miso
port 21 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 mosi
port 22 nsew
flabel metal3 s 11322 9528 12122 9648 0 FreeSans 600 0 0 0 sclk
port 23 nsew
<< properties >>
string FIXED_BBOX 0 0 12122 14266
<< end >>
